.include ../../../tech_files/TSMC_180nm.txt
.include ../../ckt_blocks/d_ff/cmos/d_ff_cmos.cir
.include ../../ckt_blocks/pg_gen/cmos/pg_gen_cmos.cir
.include ../../ckt_blocks/cla_gen/cmos/cla_gen_cmos.cir
.include ../../ckt_blocks/sum_gen/cmos/sum_gen_cmos.cir

.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={20*LAMBDA}
.param width_P={2.5*width_N}
.param length={2*LAMBDA}
.global gnd vdd

VDD vdd gnd SUPPLY
vinClk clk gnd PULSE(0 SUPPLY 10ns 1ps 1ps 10ns 20ns)
vinA3 A3 gnd PWL(0ns 0V 8ns     0V)
vinA2 A2 gnd PWL(0ns 0V 8ns     0V)
vinA1 A1 gnd PWL(0ns 0V 8ns SUPPLY)
vinA0 A0 gnd PWL(0ns 0V 8ns     0V)
vinB3 B3 gnd PWL(0ns 0V 8ns     0V)
vinB2 B2 gnd PWL(0ns 0V 8ns SUPPLY)
vinB1 B1 gnd PWL(0ns 0V 8ns     0V)
vinB0 B0 gnd PWL(0ns 0V 8ns     0V)
vinC  C  gnd PWL(0ns 0V 8ns     0V)

Xdffa3 A3 clk Q3a Q3ai d_ff_cmos
Xdffa2 A2 clk Q2a Q2ai d_ff_cmos
Xdffa1 A1 clk Q1a Q1ai d_ff_cmos
Xdffa0 A0 clk Q0a Q0ai d_ff_cmos
Xdffb3 B3 clk Q3b Q3bi d_ff_cmos
Xdffb2 B2 clk Q2b Q2bi d_ff_cmos
Xdffb1 B1 clk Q1b Q1bi d_ff_cmos
Xdffb0 B0 clk Q0b Q0bi d_ff_cmos
Xdffc   C clk  Qc  Qci d_ff_cmos

Xpg  A3 A2 A1 A0 B3 B2 B1 B0 P3 P2 P1 P0 G3 G2 G1 G0 pg_gen_cmos
Xcla  C G1 P1 G2 P2 G3 P3 C2 C3 C4 cla_gen_cmos
Xsum P3 P2 P1 P0 C3 C2 C1 C0 S3 S2 S1 S0 sum_gen_cmos

* .tran 1n 640n 

* .measure tran t_in WHEN v(A3)=0.5*SUPPLY CROSS=1
* .measure tran t_out WHEN v(G2)=0.5*SUPPLY CROSS=16
* .measure tran t_delay PARAM='t_out-t_in'

* .control
*     set hcopypscolor = 1
*     set color0=beige
*     set color1=black
*     set color2=blue
*     set color3=darkgreen
*     set color4=darkred
*     set color5=darkviolet
*     set color6=darkorange

*     run
*     plot v(A3)+30 v(A2)+28 v(A1)+26 v(A0)+24 v(B3)+22 v(B2)+20 v(B1)+18 v(B0)+16 v(P3)+14 v(P2)+12 v(P1)+10 v(P0)+8 v(G3)+6 v(G2)+4 v(G1)+2 v(G0) 
* .endc