.include ../../../../tech_files/TSMC_180nm.txt

.param SUPPLY=1.8
.global gnd vdd

VDD vdd gnd SUPPLY
vinA A gnd PULSE(0 SUPPLY 10ns 1ps 1ps 10ns 20ns)
vinB B gnd PULSE(0 SUPPLY  5ns 1ps 1ps  5ns 10ns)

.option scale=0.09u

M1000 a_7_0# B vdd w_n6_n6# CMOSP w=50 l=2
+  ad=500 pd=220 as=250 ps=110
M1001 Y A a_7_0# w_n6_n6# CMOSP w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1002 Y B gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=200 ps=100
M1003 Y A gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 A Y 0.05fF
C1 a_7_0# Y 1.03fF
C2 a_7_0# B 0.02fF
C3 a_7_0# vdd 1.03fF
C4 Y gnd 0.71fF
C5 Y w_n6_n6# 0.12fF
C6 B w_n6_n6# 0.06fF
C7 A gnd 0.05fF
C8 A w_n6_n6# 0.06fF
C9 w_n6_n6# vdd 0.12fF
C10 Y B 0.24fF
C11 a_7_0# w_n6_n6# 0.22fF
C12 gnd Gnd 0.15fF
C13 Y Gnd 0.15fF
C14 a_7_0# Gnd 0.00fF
C15 vdd Gnd 0.01fF
C16 B Gnd 0.17fF
C17 A Gnd 0.17fF
C18 w_n6_n6# Gnd 4.50fF

.tran 1n 20n 

.measure tran t_in WHEN v(B)=0.5*SUPPLY CROSS=1
.measure tran t_out WHEN v(Y)=0.5*SUPPLY CROSS=1
.measure tran t_delay PARAM='t_out-t_in'

.control
    set hcopypscolor = 1
    set color0=beige
    set color1=black
    set color2=blue
    set color3=darkgreen
    set color4=darkred
    set color5=darkviolet
    set color6=darkorange

    run
    plot v(A)+4 v(B)+2 v(Y)
    set curplottitle="2023102019"
    hardcopy nor_cmos_post_tran.eps v(A)+4 v(B)+2 v(Y)
.endc