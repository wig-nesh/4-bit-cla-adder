* SPICE3 file created from nand_5_cmos.ext - technology: scmos

.option scale=0.09u

M1000 a_39_n62# C a_23_n62# Gnd nfet w=20 l=2
+  ad=200 pd=100 as=200 ps=100
M1001 Y A vdd w_n6_n6# pfet w=50 l=2
+  ad=1250 pd=550 as=1250 ps=550
M1002 Y C vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 Y B vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_55_n62# D a_39_n62# Gnd nfet w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1005 Y E a_55_n62# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1006 Y E vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_7_n62# A gnd Gnd nfet w=20 l=2
+  ad=200 pd=100 as=100 ps=50
M1008 Y D vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_23_n62# B a_7_n62# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 A E 0.08fF
C1 Y D 0.08fF
C2 a_55_n62# a_39_n62# 0.21fF
C3 B A 0.27fF
C4 C w_n6_n6# 0.06fF
C5 a_55_n62# gnd 0.07fF
C6 C E 0.08fF
C7 B C 0.49fF
C8 Y gnd 0.03fF
C9 E a_23_n62# 0.16fF
C10 gnd a_39_n62# 0.07fF
C11 a_7_n62# a_23_n62# 0.21fF
C12 Y A 0.05fF
C13 vdd Y 4.90fF
C14 w_n6_n6# E 0.06fF
C15 A D 0.08fF
C16 Y C 0.08fF
C17 B w_n6_n6# 0.06fF
C18 B E 0.08fF
C19 C D 0.71fF
C20 a_7_n62# E 0.16fF
C21 a_23_n62# a_39_n62# 0.21fF
C22 a_55_n62# E 0.16fF
C23 gnd a_23_n62# 0.07fF
C24 vdd A 0.02fF
C25 Y w_n6_n6# 0.37fF
C26 Y E 0.13fF
C27 C A 0.08fF
C28 w_n6_n6# D 0.06fF
C29 Y B 0.26fF
C30 D E 0.93fF
C31 B D 0.08fF
C32 E a_39_n62# 0.16fF
C33 gnd E 0.05fF
C34 Y a_55_n62# 0.21fF
C35 gnd a_7_n62# 0.27fF
C36 w_n6_n6# A 0.06fF
C37 vdd w_n6_n6# 0.45fF
