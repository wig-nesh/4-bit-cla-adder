.include ../../../tech_files/TSMC_180nm.txt

.param SUPPLY=1.8
.global gnd vdd

.option scale=0.09u

.subckt inv_cmos IN w_0_0# gnd vdd OUT
M1000 OUT IN vdd w_0_0# pfet w=50 l=2
+  ad=250 pd=110 as=250 ps=110
M1001 OUT IN gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
C0 OUT gnd 0.21fF
C1 w_0_0# OUT 0.07fF
C2 vdd OUT 0.52fF
C3 IN gnd 0.05fF
C4 w_0_0# IN 0.06fF
C5 IN vdd 0.02fF
C6 w_0_0# vdd 0.07fF
C7 IN OUT 0.05fF
C8 gnd Gnd 0.06fF
C9 OUT Gnd 0.05fF
C10 vdd Gnd 0.00fF
C11 IN Gnd 0.13fF
C12 w_0_0# Gnd 1.49fF
.ends

.subckt nor_3_cmos a_23_0# Y a_7_0# gnd A B C
M1000 a_7_0# A vdd w_n6_n6# pfet w=150 l=2
+  ad=1500 pd=620 as=750 ps=310
M1001 Y C a_23_0# w_n6_n6# pfet w=150 l=2
+  ad=750 pd=310 as=1500 ps=620
M1002 a_23_0# B a_7_0# w_n6_n6# pfet w=150 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 Y A gnd Gnd nfet w=20 l=2
+  ad=300 pd=150 as=300 ps=150
M1004 Y B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 Y C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vdd a_7_0# 1.55fF
C1 a_7_0# a_23_0# 1.55fF
C2 w_n6_n6# a_7_0# 0.32fF
C3 B a_7_0# 0.02fF
C4 C a_23_0# 0.02fF
C5 w_n6_n6# C 0.06fF
C6 C Y 0.24fF
C7 w_n6_n6# A 0.06fF
C8 A Y 0.05fF
C9 A gnd 0.05fF
C10 w_n6_n6# vdd 0.17fF
C11 w_n6_n6# a_23_0# 0.32fF
C12 a_23_0# Y 1.55fF
C13 w_n6_n6# B 0.06fF
C14 w_n6_n6# Y 0.17fF
C15 B Y 0.19fF
C16 Y gnd 1.21fF
C17 gnd Gnd 0.23fF
C18 Y Gnd 0.22fF
C19 a_23_0# Gnd 0.00fF
C20 a_7_0# Gnd 0.00fF
C21 vdd Gnd 0.01fF
C22 C Gnd 0.17fF
C23 B Gnd 0.17fF
C24 A Gnd 0.17fF
C25 w_n6_n6# Gnd 9.11fF
.ends

.subckt nand_3_cmos w_n6_n6# a_7_n81# Y gnd A vdd B C a_23_n81#
M1000 Y A vdd w_n6_n6# pfet w=50 l=2
+  ad=750 pd=330 as=750 ps=330
M1001 Y C vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 Y B vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_7_n81# A gnd Gnd nfet w=60 l=2
+  ad=600 pd=260 as=300 ps=130
M1004 a_23_n81# B a_7_n81# Gnd nfet w=60 l=2
+  ad=600 pd=260 as=0 ps=0
M1005 Y C a_23_n81# Gnd nfet w=60 l=2
+  ad=300 pd=130 as=0 ps=0
C0 w_n6_n6# A 0.06fF
C1 C Y 0.24fF
C2 B a_7_n81# 0.10fF
C3 vdd Y 2.69fF
C4 A vdd 0.02fF
C5 A Y 0.05fF
C6 a_23_n81# C 0.10fF
C7 w_n6_n6# B 0.06fF
C8 w_n6_n6# C 0.06fF
C9 a_23_n81# Y 0.62fF
C10 gnd a_7_n81# 0.62fF
C11 w_n6_n6# vdd 0.25fF
C12 a_23_n81# a_7_n81# 0.62fF
C13 w_n6_n6# Y 0.22fF
C14 B Y 0.19fF
C15 a_23_n81# Gnd 0.14fF
C16 a_7_n81# Gnd 0.14fF
C17 gnd Gnd 0.10fF
C18 Y Gnd 0.20fF
C19 vdd Gnd 0.08fF
C20 C Gnd 0.17fF
C21 B Gnd 0.17fF
C22 A Gnd 0.17fF
C23 w_n6_n6# Gnd 3.49fF
.ends

.subckt nor_4_cmos Y A vdd B C D
M1000 Y D gnd Gnd nfet w=20 l=2
+  ad=400 pd=200 as=400 ps=200
M1001 a_7_0# A vdd w_n6_n6# pfet w=200 l=2
+  ad=2000 pd=820 as=1000 ps=410
M1002 a_39_0# C a_23_0# w_n6_n6# pfet w=200 l=2
+  ad=2000 pd=820 as=2000 ps=820
M1003 a_23_0# B a_7_0# w_n6_n6# pfet w=200 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 Y A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 Y B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 Y C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 Y D a_39_0# w_n6_n6# pfet w=200 l=2
+  ad=1000 pd=410 as=0 ps=0
C0 Y gnd 1.71fF
C1 w_n6_n6# B 0.06fF
C2 w_n6_n6# vdd 0.22fF
C3 a_7_0# vdd 2.06fF
C4 A gnd 0.05fF
C5 C Y 0.19fF
C6 a_23_0# w_n6_n6# 0.42fF
C7 D Y 0.24fF
C8 C w_n6_n6# 0.06fF
C9 a_23_0# a_39_0# 2.06fF
C10 a_7_0# a_23_0# 2.06fF
C11 D w_n6_n6# 0.06fF
C12 w_n6_n6# Y 0.22fF
C13 a_39_0# Y 2.06fF
C14 A Y 0.05fF
C15 a_39_0# w_n6_n6# 0.42fF
C16 B Y 0.19fF
C17 a_7_0# w_n6_n6# 0.42fF
C18 w_n6_n6# A 0.06fF
C19 gnd Gnd 0.32fF
C20 Y Gnd 0.30fF
C21 a_39_0# Gnd 0.00fF
C22 a_23_0# Gnd 0.00fF
C23 a_7_0# Gnd 0.00fF
C24 vdd Gnd 0.01fF
C25 D Gnd 0.17fF
C26 C Gnd 0.17fF
C27 B Gnd 0.17fF
C28 A Gnd 0.17fF
C29 w_n6_n6# Gnd 15.33fF
.ends

.subckt nand_cmos w_n6_n6# a_7_n61# Y A vdd B
M1000 a_7_n61# A gnd Gnd nfet w=40 l=2
+  ad=400 pd=180 as=200 ps=90
M1001 Y B a_7_n61# Gnd nfet w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1002 Y A vdd w_n6_n6# pfet w=50 l=2
+  ad=500 pd=220 as=500 ps=220
M1003 Y B vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_n6_n6# B 0.06fF
C1 vdd Y 1.60fF
C2 B Y 0.24fF
C3 a_7_n61# gnd 0.45fF
C4 w_n6_n6# Y 0.15fF
C5 A vdd 0.02fF
C6 w_n6_n6# A 0.06fF
C7 a_7_n61# B 0.05fF
C8 A Y 0.05fF
C9 a_7_n61# Y 0.41fF
C10 w_n6_n6# vdd 0.16fF
C11 a_7_n61# Gnd 0.13fF
C12 gnd Gnd 0.07fF
C13 Y Gnd 0.14fF
C14 vdd Gnd 0.05fF
C15 B Gnd 0.17fF
C16 A Gnd 0.17fF
C17 w_n6_n6# Gnd 2.49fF
.ends

.subckt nor_cmos Y a_7_0# A B
M1000 a_7_0# A vdd w_n6_n6# pfet w=100 l=2
+  ad=1000 pd=420 as=500 ps=210
M1001 Y B a_7_0# w_n6_n6# pfet w=100 l=2
+  ad=500 pd=210 as=0 ps=0
M1002 Y A gnd Gnd nfet w=20 l=2
+  ad=200 pd=100 as=200 ps=100
M1003 Y B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 vdd w_n6_n6# 0.12fF
C1 Y B 0.24fF
C2 Y A 0.05fF
C3 a_7_0# w_n6_n6# 0.22fF
C4 Y a_7_0# 1.03fF
C5 Y gnd 0.71fF
C6 B a_7_0# 0.02fF
C7 gnd A 0.05fF
C8 Y w_n6_n6# 0.12fF
C9 vdd a_7_0# 1.03fF
C10 B w_n6_n6# 0.06fF
C11 w_n6_n6# A 0.06fF
C12 gnd Gnd 0.15fF
C13 Y Gnd 0.15fF
C14 a_7_0# Gnd 0.00fF
C15 vdd Gnd 0.01fF
C16 B Gnd 0.17fF
C17 A Gnd 0.17fF
C18 w_n6_n6# Gnd 4.50fF
.ends

.subckt nand_4_cmos w_n6_n6# a_7_n101# a_7_0# A vdd a_39_n101# B a_23_n101# C D
M1000 a_7_0# D a_39_n101# Gnd nfet w=80 l=2
+  ad=400 pd=170 as=800 ps=340
M1001 a_7_0# A vdd w_n6_n6# pfet w=50 l=2
+  ad=1000 pd=440 as=1000 ps=440
M1002 a_7_0# C vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_7_0# B vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_7_n101# A gnd Gnd nfet w=80 l=2
+  ad=800 pd=340 as=400 ps=170
M1005 a_39_n101# C a_23_n101# Gnd nfet w=80 l=2
+  ad=0 pd=0 as=800 ps=340
M1006 a_23_n101# B a_7_n101# Gnd nfet w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_7_0# D vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
C0 C a_23_n101# 0.10fF
C1 a_23_n101# a_39_n101# 0.82fF
C2 D a_39_n101# 0.10fF
C3 gnd a_7_n101# 0.82fF
C4 vdd a_7_0# 3.78fF
C5 vdd w_n6_n6# 0.34fF
C6 B a_7_0# 0.19fF
C7 B w_n6_n6# 0.06fF
C8 a_7_n101# a_23_n101# 0.82fF
C9 vdd A 0.02fF
C10 w_n6_n6# a_7_0# 0.29fF
C11 A a_7_0# 0.05fF
C12 w_n6_n6# A 0.06fF
C13 C a_7_0# 0.19fF
C14 C w_n6_n6# 0.06fF
C15 D a_7_0# 0.24fF
C16 B a_7_n101# 0.10fF
C17 D w_n6_n6# 0.06fF
C18 a_7_0# a_39_n101# 0.82fF
C19 a_39_n101# Gnd 0.18fF
C20 a_23_n101# Gnd 0.18fF
C21 a_7_n101# Gnd 0.18fF
C22 gnd Gnd 0.12fF
C23 a_7_0# Gnd 0.02fF
C24 vdd Gnd 0.03fF
C25 D Gnd 0.17fF
C26 C Gnd 0.15fF
C27 B Gnd 0.15fF
C28 A Gnd -0.00fF
C29 w_n6_n6# Gnd 4.48fF
.ends

.subckt nor_5_cmos a_23_0# w_n6_n6# Y a_7_0# A vdd B C D a_39_0# E a_55_0#
M1000 a_7_0# A vdd w_n6_n6# pfet w=250 l=2
+  ad=2500 pd=1020 as=1250 ps=510
M1001 a_39_0# C a_23_0# w_n6_n6# pfet w=250 l=2
+  ad=2500 pd=1020 as=2500 ps=1020
M1002 a_23_0# B a_7_0# w_n6_n6# pfet w=250 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 Y D gnd Gnd nfet w=20 l=2
+  ad=500 pd=250 as=500 ps=250
M1004 Y E gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 Y A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 Y E a_55_0# w_n6_n6# pfet w=250 l=2
+  ad=1250 pd=510 as=2500 ps=1020
M1007 Y B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 a_55_0# D a_39_0# w_n6_n6# pfet w=250 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 Y C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_n6_n6# E 0.06fF
C1 Y C 0.19fF
C2 a_39_0# D 0.02fF
C3 Y D 0.19fF
C4 w_n6_n6# B 0.06fF
C5 Y E 0.24fF
C6 a_55_0# w_n6_n6# 0.52fF
C7 Y B 0.19fF
C8 A gnd 0.05fF
C9 a_7_0# w_n6_n6# 0.52fF
C10 a_55_0# a_39_0# 2.58fF
C11 a_7_0# a_23_0# 2.58fF
C12 Y gnd 2.21fF
C13 a_55_0# Y 2.58fF
C14 a_7_0# vdd 2.58fF
C15 a_23_0# w_n6_n6# 0.52fF
C16 a_55_0# E 0.02fF
C17 w_n6_n6# A 0.06fF
C18 a_39_0# w_n6_n6# 0.52fF
C19 a_23_0# a_39_0# 2.58fF
C20 vdd w_n6_n6# 0.27fF
C21 w_n6_n6# C 0.06fF
C22 a_23_0# C 0.02fF
C23 Y w_n6_n6# 0.27fF
C24 w_n6_n6# D 0.06fF
C25 Y A 0.05fF
C26 a_7_0# B 0.02fF
C27 gnd Gnd 0.41fF
C28 Y Gnd 0.38fF
C29 a_55_0# Gnd -0.00fF
C30 a_39_0# Gnd -0.00fF
C31 a_23_0# Gnd -0.00fF
C32 a_7_0# Gnd -0.00fF
C33 vdd Gnd 0.01fF
C34 E Gnd 0.17fF
C35 D Gnd 0.17fF
C36 C Gnd 0.17fF
C37 B Gnd 0.17fF
C38 A Gnd 0.17fF
C39 w_n6_n6# Gnd 23.16fF
.ends

.subckt nand_5_cmos a_7_n121# w_n6_n6# a_55_n121# Y gnd a_39_n121# a_23_n121# A vdd
+ B C D E
M1000 Y A vdd w_n6_n6# pfet w=50 l=2
+  ad=1250 pd=550 as=1250 ps=550
M1001 Y C vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 Y B vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 Y E a_55_n121# Gnd nfet w=100 l=2
+  ad=500 pd=210 as=1000 ps=420
M1004 a_55_n121# D a_39_n121# Gnd nfet w=100 l=2
+  ad=0 pd=0 as=1000 ps=420
M1005 Y E vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 Y D vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_7_n121# A gnd Gnd nfet w=100 l=2
+  ad=1000 pd=420 as=500 ps=210
M1008 a_39_n121# C a_23_n121# Gnd nfet w=100 l=2
+  ad=0 pd=0 as=1000 ps=420
M1009 a_23_n121# B a_7_n121# Gnd nfet w=100 l=2
+  ad=0 pd=0 as=0 ps=0
C0 C a_23_n121# 0.10fF
C1 a_39_n121# a_55_n121# 1.03fF
C2 a_23_n121# a_39_n121# 1.03fF
C3 Y w_n6_n6# 0.37fF
C4 w_n6_n6# D 0.06fF
C5 B w_n6_n6# 0.06fF
C6 Y a_55_n121# 1.03fF
C7 Y E 0.24fF
C8 Y A 0.05fF
C9 B a_7_n121# 0.10fF
C10 Y vdd 4.87fF
C11 C Y 0.19fF
C12 a_39_n121# D 0.10fF
C13 w_n6_n6# E 0.06fF
C14 gnd a_7_n121# 1.03fF
C15 w_n6_n6# A 0.06fF
C16 E a_55_n121# 0.10fF
C17 vdd w_n6_n6# 0.42fF
C18 C w_n6_n6# 0.06fF
C19 a_7_n121# a_23_n121# 1.03fF
C20 vdd A 0.02fF
C21 Y D 0.19fF
C22 B Y 0.19fF
C23 a_55_n121# Gnd 0.22fF
C24 a_39_n121# Gnd 0.22fF
C25 a_23_n121# Gnd 0.22fF
C26 a_7_n121# Gnd 0.22fF
C27 gnd Gnd 0.14fF
C28 Y Gnd 0.28fF
C29 vdd Gnd 0.14fF
C30 E Gnd 0.13fF
C31 D Gnd 0.13fF
C32 C Gnd 0.13fF
C33 B Gnd 0.13fF
C34 A Gnd 0.13fF
C35 w_n6_n6# Gnd 5.48fF
.ends

.subckt cla_gen_cmos_unrouted
Xinv_cmos_3 nand_cmos_0/Y inv_cmos_3/w_0_0# inv_cmos_3/gnd inv_cmos_3/vdd d inv_cmos
Xinv_cmos_4 inv_cmos_4/IN inv_cmos_4/w_0_0# inv_cmos_4/gnd inv_cmos_4/vdd e inv_cmos
Xinv_cmos_6 nand_cmos_1/Y inv_cmos_6/w_0_0# inv_cmos_6/gnd inv_cmos_6/vdd g inv_cmos
Xinv_cmos_5 inv_cmos_5/IN inv_cmos_5/w_0_0# inv_cmos_5/gnd inv_cmos_5/vdd f inv_cmos
Xinv_cmos_7 inv_cmos_7/IN inv_cmos_7/w_0_0# inv_cmos_7/gnd inv_cmos_7/vdd h inv_cmos
Xnor_3_cmos_0 nor_3_cmos_0/a_23_0# m nor_3_cmos_0/a_7_0# nor_3_cmos_0/gnd h i G1 nor_3_cmos
Xinv_cmos_8 nand_cmos_2/Y inv_cmos_8/w_0_0# inv_cmos_8/gnd inv_cmos_8/vdd i inv_cmos
Xinv_cmos_9 nand_cmos_3/Y inv_cmos_9/w_0_0# inv_cmos_9/gnd inv_cmos_9/vdd j inv_cmos
Xnand_3_cmos_0 inv_cmos_2/w_0_0# nand_3_cmos_0/a_7_n81# inv_cmos_2/IN nand_3_cmos_0/gnd
+ P3 nand_3_cmos_0/vdd P2 G1 nand_3_cmos_0/a_23_n81# nand_3_cmos
Xnor_4_cmos_0 l e nor_4_cmos_0/vdd f g G2 nor_4_cmos
Xnand_3_cmos_1 inv_cmos_5/w_0_0# nand_3_cmos_1/a_7_n81# inv_cmos_5/IN nand_3_cmos_1/gnd
+ P2 nand_3_cmos_1/vdd P1 G0 nand_3_cmos_1/a_23_n81# nand_3_cmos
Xnand_3_cmos_2 inv_cmos_7/w_0_0# nand_3_cmos_2/a_7_n81# inv_cmos_7/IN nand_5_cmos_0/gnd
+ P1 nand_3_cmos_2/vdd P0 C0 nand_3_cmos_2/a_23_n81# nand_3_cmos
Xnand_cmos_1 inv_cmos_6/w_0_0# nand_cmos_1/a_7_n61# nand_cmos_1/Y P2 nand_cmos_1/vdd
+ G1 nand_cmos
Xnand_cmos_0 inv_cmos_3/w_0_0# nand_cmos_0/a_7_n61# nand_cmos_0/Y P3 nand_cmos_0/vdd
+ G2 nand_cmos
Xnand_cmos_2 inv_cmos_8/w_0_0# nand_cmos_2/a_7_n61# nand_cmos_2/Y P1 nand_cmos_2/vdd
+ G0 nand_cmos
Xinv_cmos_11 l inv_cmos_11/w_0_0# inv_cmos_11/gnd inv_cmos_11/vdd C3 inv_cmos
Xinv_cmos_10 k inv_cmos_10/w_0_0# inv_cmos_10/gnd inv_cmos_10/vdd C4 inv_cmos
Xnor_cmos_0 n nor_cmos_0/a_7_0# j G0 nor_cmos
Xnand_4_cmos_0 inv_cmos_1/w_0_0# nand_4_cmos_0/a_7_n101# inv_cmos_1/IN P3 nand_4_cmos_0/vdd
+ nand_4_cmos_0/a_39_n101# P2 nand_4_cmos_0/a_23_n101# P1 G0 nand_4_cmos
Xnand_cmos_3 inv_cmos_9/w_0_0# nand_cmos_3/a_7_n61# nand_cmos_3/Y P0 nand_cmos_3/vdd
+ C0 nand_cmos
Xnand_4_cmos_1 inv_cmos_4/w_0_0# nand_4_cmos_1/a_7_n101# inv_cmos_4/IN P2 nand_4_cmos_1/vdd
+ nand_4_cmos_1/a_39_n101# P1 nand_4_cmos_1/a_23_n101# P0 C0 nand_4_cmos
Xinv_cmos_12 m inv_cmos_12/w_0_0# inv_cmos_12/gnd inv_cmos_12/vdd C2 inv_cmos
Xnor_5_cmos_0 nor_5_cmos_0/a_23_0# nor_5_cmos_0/w_n6_n6# k nor_5_cmos_0/a_7_0# a nor_5_cmos_0/vdd
+ b c d nor_5_cmos_0/a_39_0# G3 nor_5_cmos_0/a_55_0# nor_5_cmos
Xinv_cmos_13 n inv_cmos_13/w_0_0# inv_cmos_13/gnd inv_cmos_13/vdd C1 inv_cmos
Xnand_5_cmos_0 nand_5_cmos_0/a_7_n121# inv_cmos_0/w_0_0# nand_5_cmos_0/a_55_n121#
+ inv_cmos_0/IN nand_5_cmos_0/gnd nand_5_cmos_0/a_39_n121# nand_5_cmos_0/a_23_n121#
+ P3 nand_5_cmos_0/vdd P2 P1 P0 C0 nand_5_cmos
Xinv_cmos_0 inv_cmos_0/IN inv_cmos_0/w_0_0# inv_cmos_0/gnd inv_cmos_0/vdd a inv_cmos
Xinv_cmos_1 inv_cmos_1/IN inv_cmos_1/w_0_0# inv_cmos_1/gnd inv_cmos_1/vdd b inv_cmos
Xinv_cmos_2 inv_cmos_2/IN inv_cmos_2/w_0_0# inv_cmos_2/gnd inv_cmos_2/vdd c inv_cmos
C0 nand_3_cmos_1/vdd nand_4_cmos_0/vdd 0.21fF
C1 a P3 0.02fF
C2 G0 nand_cmos_2/a_7_n61# 0.05fF
C3 G1 nand_cmos_1/Y 0.05fF
C4 e P2 0.02fF
C5 nand_3_cmos_1/a_23_n81# G0 0.05fF
C6 P1 P2 0.08fF
C7 nand_cmos_0/Y inv_cmos_3/gnd 0.30fF
C8 C0 inv_cmos_0/IN 0.05fF
C9 inv_cmos_9/vdd nand_cmos_3/Y 0.52fF
C10 C4 m 0.02fF
C11 nor_3_cmos_0/a_7_0# i 0.02fF
C12 inv_cmos_4/IN inv_cmos_4/w_0_0# 0.00fF
C13 d k 0.05fF
C14 G3 nor_5_cmos_0/a_55_0# 0.02fF
C15 P1 inv_cmos_1/IN 0.05fF
C16 G0 nand_4_cmos_0/a_39_n101# 0.05fF
C17 P1 P0 0.08fF
C18 nand_3_cmos_0/vdd nor_4_cmos_0/vdd 0.04fF
C19 G1 inv_cmos_2/IN 0.05fF
C20 nor_3_cmos_0/gnd nand_3_cmos_0/a_7_n81# 0.01fF
C21 nand_cmos_2/Y G0 0.05fF
C22 P1 inv_cmos_0/IN 0.05fF
C23 inv_cmos_4/IN P0 0.05fF
C24 C0 nand_5_cmos_0/a_55_n121# 0.05fF
C25 C0 nand_4_cmos_1/a_39_n101# 0.05fF
C26 inv_cmos_6/gnd nand_cmos_1/Y 0.30fF
C27 inv_cmos_6/vdd nand_cmos_1/Y 0.52fF
C28 G1 i 0.04fF
C29 nor_5_cmos_0/w_n6_n6# nor_5_cmos_0/vdd -0.00fF
C30 b k 0.05fF
C31 d nor_5_cmos_0/a_39_0# 0.02fF
C32 nand_4_cmos_1/vdd nand_5_cmos_0/vdd 0.54fF
C33 nor_3_cmos_0/gnd inv_cmos_2/IN 0.02fF
C34 nand_cmos_2/Y inv_cmos_8/w_0_0# -0.00fF
C35 nand_cmos_0/Y G2 0.05fF
C36 nand_4_cmos_0/a_7_n101# P2 0.05fF
C37 nand_3_cmos_1/a_7_n81# P1 0.05fF
C38 inv_cmos_5/gnd inv_cmos_5/IN 0.30fF
C39 nand_cmos_2/Y inv_cmos_8/gnd 0.30fF
C40 P0 nand_5_cmos_0/a_39_n121# 0.05fF
C41 P0 nand_4_cmos_1/a_23_n101# 0.05fF
C42 G1 m 0.05fF
C43 C2 n 0.02fF
C44 C0 nand_cmos_3/a_7_n61# 0.05fF
C45 inv_cmos_1/IN inv_cmos_1/gnd 0.30fF
C46 P2 nand_5_cmos_0/a_7_n121# 0.05fF
C47 c nor_5_cmos_0/a_23_0# 0.02fF
C48 P1 nand_4_cmos_0/a_23_n101# 0.05fF
C49 G0 inv_cmos_1/IN 0.05fF
C50 G1 nand_3_cmos_0/a_23_n81# 0.05fF
C51 b P3 0.02fF
C52 G0 nor_cmos_0/a_7_0# 0.02fF
C53 inv_cmos_1/IN P2 0.05fF
C54 inv_cmos_5/IN P1 0.05fF
C55 inv_cmos_5/vdd inv_cmos_5/IN 0.52fF
C56 nand_cmos_2/Y inv_cmos_8/vdd 0.52fF
C57 f P2 0.02fF
C58 P1 nand_5_cmos_0/a_23_n121# 0.05fF
C59 P1 nand_4_cmos_1/a_7_n101# 0.05fF
C60 nand_cmos_1/vdd inv_cmos_1/vdd 0.04fF
C61 C0 nand_cmos_3/Y 0.05fF
C62 inv_cmos_1/IN inv_cmos_1/vdd 0.52fF
C63 inv_cmos_4/vdd nand_5_cmos_0/vdd 0.04fF
C64 inv_cmos_4/vdd inv_cmos_4/IN 0.52fF
C65 P2 inv_cmos_0/IN 0.05fF
C66 b nor_5_cmos_0/a_7_0# 0.02fF
C67 d G3 0.04fF
C68 inv_cmos_7/IN P0 0.05fF
C69 G3 k 0.05fF
C70 G1 P2 0.04fF
C71 C0 nand_3_cmos_2/a_23_n81# 0.07fF
C72 nor_3_cmos_0/gnd nand_3_cmos_0/a_23_n81# 0.05fF
C73 P0 inv_cmos_0/IN 0.05fF
C74 inv_cmos_4/IN C0 0.05fF
C75 inv_cmos_0/IN inv_cmos_0/gnd 0.30fF
C76 g f 0.04fF
C77 inv_cmos_1/IN inv_cmos_1/w_0_0# 0.00fF
C78 G0 n 0.05fF
C79 c d 0.04fF
C80 inv_cmos_7/IN inv_cmos_7/w_0_0# -0.00fF
C81 c k 0.05fF
C82 inv_cmos_5/w_0_0# inv_cmos_5/IN 0.00fF
C83 G2 nand_cmos_0/a_7_n61# 0.04fF
C84 inv_cmos_5/vdd nand_4_cmos_0/vdd 0.04fF
C85 inv_cmos_2/IN inv_cmos_2/gnd 0.30fF
C86 P0 nand_3_cmos_2/a_7_n81# 0.07fF
C87 inv_cmos_5/IN G0 0.05fF
C88 nand_cmos_0/Y inv_cmos_3/vdd 0.52fF
C89 inv_cmos_4/IN P1 0.05fF
C90 inv_cmos_7/IN inv_cmos_7/gnd 0.30fF
C91 inv_cmos_0/IN inv_cmos_0/vdd 0.52fF
C92 f l 0.05fF
C93 b c 0.04fF
C94 g G2 0.04fF
C95 nand_3_cmos_0/a_7_n81# P2 0.05fF
C96 g l 0.05fF
C97 inv_cmos_2/IN inv_cmos_2/vdd 0.52fF
C98 inv_cmos_4/gnd inv_cmos_4/IN 0.30fF
C99 c P3 0.02fF
C100 G1 nand_cmos_1/a_7_n61# 0.04fF
C101 i m 0.05fF
C102 inv_cmos_7/IN inv_cmos_7/vdd 0.52fF
C103 inv_cmos_9/gnd nand_cmos_3/Y 0.30fF
C104 inv_cmos_6/vdd nand_3_cmos_0/vdd 0.04fF
C105 inv_cmos_7/IN C0 0.05fF
C106 l G2 0.05fF
C107 inv_cmos_2/IN P2 0.05fF
C108 G1 nor_3_cmos_0/a_23_0# 0.02fF
C109 inv_cmos_2/IN inv_cmos_2/w_0_0# 0.00fF
C110 P0 C0 0.12fF
C111 P1 G0 0.08fF
C112 inv_cmos_0/IN Gnd 0.01fF
C113 P2 Gnd 0.02fF
C114 P3 Gnd 0.06fF
C115 C1 Gnd 0.02fF
C116 n Gnd 0.00fF
C117 k Gnd 0.04fF
C118 G3 Gnd -0.01fF
C119 d Gnd -0.01fF
C120 c Gnd 0.04fF
C121 b Gnd -0.06fF
C122 a Gnd 0.02fF
C123 C2 Gnd 0.02fF
C124 m Gnd 0.04fF
C125 nand_cmos_3/Y Gnd 0.00fF
C126 inv_cmos_1/IN Gnd 0.01fF
C127 C4 Gnd 0.02fF
C128 C3 Gnd 0.02fF
C129 G0 Gnd -0.04fF
C130 G2 Gnd 0.00fF
C131 nand_cmos_1/Y Gnd -0.02fF
C132 C0 Gnd -0.01fF
C133 P0 Gnd 0.05fF
C134 P1 Gnd 0.13fF
C135 inv_cmos_5/IN Gnd 0.01fF
C136 l Gnd 0.04fF
C137 inv_cmos_2/IN Gnd 0.01fF
C138 j Gnd 0.04fF
C139 i Gnd 0.04fF
C140 nand_cmos_2/Y Gnd 0.01fF
C141 G1 Gnd 0.06fF
C142 h Gnd 0.04fF
C143 inv_cmos_7/IN Gnd 0.01fF
C144 f Gnd 0.04fF
C145 g Gnd 0.04fF
C146 e Gnd 0.04fF
C147 inv_cmos_4/IN Gnd 0.01fF
C148 nand_cmos_0/Y Gnd 0.01fF
.ends

.subckt xor_optimized Y w_26_37# A B inv_cmos_0/vdd
Xinv_cmos_0 B w_26_37# inv_cmos_0/gnd inv_cmos_0/vdd inv_cmos_0/OUT inv_cmos
M1000 Y A inv_cmos_0/OUT Gnd nfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1001 Y A B w_26_37# pfet w=50 l=2
+  ad=250 pd=110 as=320 ps=110
C0 Y w_26_37# 0.07fF
C1 B inv_cmos_0/OUT 0.70fF
C2 Y inv_cmos_0/OUT 0.28fF
C3 B A 0.05fF
C4 A w_26_37# 0.10fF
C5 Y B 0.56fF
C6 B w_26_37# 0.28fF
C7 Y Gnd 0.05fF
C8 A Gnd 0.01fF
C9 inv_cmos_0/OUT Gnd 0.06fF
C10 B Gnd 0.32fF
C11 w_26_37# Gnd 1.12fF
.ends

.subckt pg_gen_optimized_unrouted
Xinv_cmos_3 nand_cmos_3/Y inv_cmos_3/w_0_0# inv_cmos_3/gnd inv_cmos_3/vdd G0 inv_cmos
Xnand_cmos_1 inv_cmos_1/w_0_0# nand_cmos_1/a_7_n61# nand_cmos_1/Y B2 inv_cmos_1/vdd
+ A2 nand_cmos
Xnand_cmos_0 inv_cmos_0/w_0_0# nand_cmos_0/a_7_n61# nand_cmos_0/Y B3 inv_cmos_0/vdd
+ A3 nand_cmos
Xnand_cmos_2 inv_cmos_2/w_0_0# nand_cmos_2/a_7_n61# nand_cmos_2/Y B1 inv_cmos_2/vdd
+ A1 nand_cmos
Xnand_cmos_3 inv_cmos_3/w_0_0# nand_cmos_3/a_7_n61# nand_cmos_3/Y B0 inv_cmos_3/vdd
+ A0 nand_cmos
Xxor_optimized_0 P3 xor_optimized_0/w_26_37# A3 B3 inv_cmos_0/vdd xor_optimized
Xxor_optimized_1 P2 xor_optimized_1/w_26_37# A2 B2 inv_cmos_1/vdd xor_optimized
Xxor_optimized_2 P1 xor_optimized_2/w_26_37# A1 B1 inv_cmos_2/vdd xor_optimized
Xxor_optimized_3 P0 xor_optimized_3/w_26_37# A0 B0 inv_cmos_3/vdd xor_optimized
Xinv_cmos_0 nand_cmos_0/Y inv_cmos_0/w_0_0# inv_cmos_0/gnd inv_cmos_0/vdd G3 inv_cmos
Xinv_cmos_1 nand_cmos_1/Y inv_cmos_1/w_0_0# inv_cmos_1/gnd inv_cmos_1/vdd G2 inv_cmos
Xinv_cmos_2 nand_cmos_2/Y inv_cmos_2/w_0_0# inv_cmos_2/gnd inv_cmos_2/vdd G1 inv_cmos
C0 inv_cmos_1/vdd nand_cmos_1/Y 0.55fF
C1 inv_cmos_1/vdd inv_cmos_1/w_0_0# 0.01fF
C2 inv_cmos_3/gnd nand_cmos_3/Y 0.30fF
C3 G2 B1 0.02fF
C4 A2 nand_cmos_1/a_7_n61# 0.04fF
C5 inv_cmos_2/vdd A1 0.16fF
C6 nand_cmos_0/Y A3 0.05fF
C7 G3 B2 0.02fF
C8 xor_optimized_1/w_26_37# A2 0.01fF
C9 inv_cmos_0/vdd inv_cmos_0/w_0_0# 0.01fF
C10 A1 xor_optimized_2/w_26_37# 0.01fF
C11 inv_cmos_1/vdd A2 0.16fF
C12 G1 B0 0.02fF
C13 nand_cmos_3/Y inv_cmos_3/vdd 0.55fF
C14 nand_cmos_3/Y A0 0.05fF
C15 nand_cmos_3/Y inv_cmos_3/w_0_0# -0.00fF
C16 A2 nand_cmos_1/Y 0.05fF
C17 nand_cmos_3/a_7_n61# A0 0.04fF
C18 nand_cmos_2/a_7_n61# A1 0.04fF
C19 nand_cmos_0/a_7_n61# A3 0.04fF
C20 nand_cmos_2/Y inv_cmos_2/gnd 0.30fF
C21 inv_cmos_0/vdd A3 0.16fF
C22 nand_cmos_2/Y inv_cmos_2/w_0_0# -0.00fF
C23 inv_cmos_0/vdd nand_cmos_0/Y 0.55fF
C24 nand_cmos_1/Y inv_cmos_1/gnd 0.30fF
C25 A3 xor_optimized_0/w_26_37# 0.01fF
C26 xor_optimized_3/w_26_37# A0 0.01fF
C27 inv_cmos_3/vdd A0 0.16fF
C28 nand_cmos_2/Y A1 0.05fF
C29 inv_cmos_3/w_0_0# inv_cmos_3/vdd 0.01fF
C30 inv_cmos_2/w_0_0# inv_cmos_2/vdd 0.01fF
C31 inv_cmos_0/w_0_0# nand_cmos_0/Y -0.00fF
C32 nand_cmos_0/Y inv_cmos_0/gnd 0.30fF
C33 nand_cmos_2/Y inv_cmos_2/vdd 0.55fF
C34 inv_cmos_3/vdd Gnd -0.31fF
C35 inv_cmos_2/vdd Gnd -0.11fF
C36 inv_cmos_1/vdd Gnd -0.14fF
C37 G1 Gnd 0.02fF
C38 G2 Gnd 0.02fF
C39 G3 Gnd 0.02fF
C40 P0 Gnd 0.02fF
C41 A0 Gnd 0.03fF
C42 B0 Gnd 0.00fF
C43 P1 Gnd 0.02fF
C44 A1 Gnd 0.03fF
C45 B1 Gnd 0.04fF
C46 P2 Gnd 0.02fF
C47 A2 Gnd 0.03fF
C48 B2 Gnd 0.04fF
C49 P3 Gnd 0.02fF
C50 A3 Gnd 0.03fF
C51 inv_cmos_0/vdd Gnd -0.11fF
C52 B3 Gnd 0.04fF
C53 nand_cmos_3/Y Gnd 0.01fF
C54 nand_cmos_2/Y Gnd 0.01fF
C55 nand_cmos_0/Y Gnd 0.01fF
C56 nand_cmos_1/Y Gnd 0.01fF
C57 G0 Gnd 0.02fF
.ends

.subckt sum_gen_optimized_unrouted
Xxor_optimized_0 S2 xor_optimized_0/w_26_37# C2 P2 xor_optimized_2/inv_cmos_0/vdd
+ xor_optimized
Xxor_optimized_1 S1 xor_optimized_1/w_26_37# C1 P1 xor_optimized_3/inv_cmos_0/vdd
+ xor_optimized
Xxor_optimized_2 S0 xor_optimized_2/w_26_37# C0 P0 xor_optimized_2/inv_cmos_0/vdd
+ xor_optimized
Xxor_optimized_3 S3 xor_optimized_3/w_26_37# C3 P3 xor_optimized_3/inv_cmos_0/vdd
+ xor_optimized
C0 P1 S2 0.08fF
C1 S0 P3 0.08fF
C2 C1 C3 0.15fF
C3 xor_optimized_0/w_26_37# C2 0.01fF
C4 xor_optimized_3/w_26_37# C3 0.01fF
C5 C0 C2 0.15fF
C6 xor_optimized_2/w_26_37# C0 0.01fF
C7 xor_optimized_1/w_26_37# C1 0.01fF
C8 S3 Gnd -0.06fF
C9 C3 Gnd -0.20fF
C10 P3 Gnd 0.02fF
C11 S0 Gnd 0.02fF
C12 C0 Gnd -0.04fF
C13 P0 Gnd 0.02fF
C14 S1 Gnd -0.06fF
C15 C1 Gnd -0.15fF
C16 P1 Gnd 0.02fF
C17 S2 Gnd 0.02fF
C18 C2 Gnd 0.01fF
C19 P2 Gnd 0.02fF
.ends

.tran 1n 6n 

.measure tran delay_S3_r TRIG V(A3) VAL=0.5*SUPPLY RISE=1 TARG V(S3) VAL=0.5*SUPPLY RISE=1
.measure tran delay_S2_r TRIG V(A2) VAL=0.5*SUPPLY RISE=1 TARG V(S2) VAL=0.5*SUPPLY RISE=1
.measure tran delay_S1_r TRIG V(A1) VAL=0.5*SUPPLY RISE=1 TARG V(S1) VAL=0.5*SUPPLY RISE=1
.measure tran delay_S0_r TRIG V(A0) VAL=0.5*SUPPLY RISE=1 TARG V(S0) VAL=0.5*SUPPLY RISE=1
.measure tran delay_C4_r TRIG V(C0) VAL=0.5*SUPPLY RISE=1 TARG V(C4) VAL=0.5*SUPPLY RISE=1
.measure tran delay_S3_f TRIG V(A3) VAL=0.5*SUPPLY FALL=1 TARG V(S3) VAL=0.5*SUPPLY FALL=1
.measure tran delay_S2_f TRIG V(A2) VAL=0.5*SUPPLY FALL=1 TARG V(S2) VAL=0.5*SUPPLY FALL=1
.measure tran delay_S1_f TRIG V(A1) VAL=0.5*SUPPLY FALL=1 TARG V(S1) VAL=0.5*SUPPLY FALL=1
.measure tran delay_S0_f TRIG V(A0) VAL=0.5*SUPPLY FALL=1 TARG V(S0) VAL=0.5*SUPPLY FALL=1
.measure tran delay_C4_f TRIG V(C0) VAL=0.5*SUPPLY FALL=1 TARG V(C4) VAL=0.5*SUPPLY FALL=1


.control
    set hcopypscolor = 1
    set color0=beige
    set color1=black
    set color2=blue
    set color3=darkgreen
    set color4=darkred
    set color5=darkviolet
    set color6=darkorange

    run
    plot v(clk)+28 v(A3)+26 v(A2)+24 v(A1)+22 v(A0)+20 v(B3)+18 v(B2)+16 v(B1)+14 v(B0)+12 v(C0)+10 v(Q3s)+8 v(S3)+8 v(Q2s)+6 v(S2)+6 v(Q1s)+4 v(S1)+4 v(Q0s)+2 v(S0)+2 v(Qco) v(C4)
    * plot v(clk)+28 v(A3)+26 v(A2)+24 v(A1)+22 v(A0)+20 v(B3)+18 v(B2)+16 v(B1)+14 v(B0)+12 v(C0)+10 v(S3)+8 v(S2)+6 v(S1)+4 v(S0)+2 v(C4)
    * plot v(clk)+28 v(A3)+26 v(A2)+24 v(A1)+22 v(A0)+20 v(B3)+18 v(B2)+16 v(B1)+14 v(B0)+12 v(C0)+10 v(Q3a)+8 v(Q2a)+6 v(Q1a)+4 v(Q0a)+2 v(Q3b) v(Q2b)-2 v(Q1b)-4 v(Q0b)-6 v(Qc0)-8
    * plot v(clk)+28 v(A3)+26 v(A2)+24 v(A1)+22 v(A0)+20 v(B3)+18 v(B2)+16 v(B1)+14 v(B0)+12 v(C0)+10 v(P3)+8 v(P2)+6 v(P1)+4 v(P0)+2 v(G3) v(G2)-2 v(G1)-4 v(G0)-6
    * plot v(clk)+28 v(A3)+26 v(A2)+24 v(A1)+22 v(A0)+20 v(B3)+18 v(B2)+16 v(B1)+14 v(B0)+12 v(C0)+10 v(C4)+8 v(C3)+6 v(C2)+4 v(C1)+2
    * plot v(clk)+28 v(A3)+26 v(A2)+24 v(A1)+22 v(A0)+20 v(B3)+18 v(B2)+16 v(B1)+14 v(B0)+12 v(C0)+10 v(S3)+8 v(S2)+6 v(S1)+4 v(S0)+2 v(C4)
.endc