.include ../../../../tech_files/TSMC_180nm.txt

.param SUPPLY=1.8
.global gnd vdd

VDD vdd gnd SUPPLY
vinA A gnd PULSE(0 SUPPLY  10ns 1ps 1ps  10ns 20ns)
vinB B gnd PULSE(0 SUPPLY   5ns 1ps 1ps   5ns 10ns)
vinC C gnd PULSE(0 SUPPLY 2.5ns 1ps 1ps 2.5ns  5ns)

.option scale=0.09u

M1000 Y A vdd w_n6_n6# CMOSP w=50 l=2
+  ad=750 pd=330 as=750 ps=330
M1001 Y C vdd w_n6_n6# CMOSP w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 Y B vdd w_n6_n6# CMOSP w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_7_n81# A gnd Gnd CMOSN w=60 l=2
+  ad=600 pd=260 as=300 ps=130
M1004 a_23_n81# B a_7_n81# Gnd CMOSN w=60 l=2
+  ad=600 pd=260 as=0 ps=0
M1005 Y C a_23_n81# Gnd CMOSN w=60 l=2
+  ad=300 pd=130 as=0 ps=0
C0 a_7_n81# a_23_n81# 0.62fF
C1 vdd Y 2.69fF
C2 B a_7_n81# 0.10fF
C3 A Y 0.05fF
C4 w_n6_n6# vdd 0.25fF
C5 w_n6_n6# A 0.06fF
C6 C a_23_n81# 0.10fF
C7 C Y 0.24fF
C8 A vdd 0.02fF
C9 w_n6_n6# C 0.06fF
C10 Y a_23_n81# 0.62fF
C11 gnd a_7_n81# 0.62fF
C12 B Y 0.19fF
C13 w_n6_n6# Y 0.22fF
C14 w_n6_n6# B 0.06fF



.tran 1n 20n 

.control
    set hcopypscolor = 1
    set color0=beige
    set color1=black
    set color2=blue
    set color3=darkgreen
    set color4=darkred
    set color5=darkviolet
    set color6=darkorange

    run
    plot v(A)+4 v(B)+2 v(C) v(Y)-2
.endc