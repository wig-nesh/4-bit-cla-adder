* SPICE3 file created from nor_3_cmos.ext - technology: scmos

.option scale=0.09u

M1000 a_7_0# A vdd w_n6_n6# pfet w=150 l=2
+  ad=1500 pd=620 as=750 ps=310
M1001 Y C a_23_0# w_n6_n6# pfet w=150 l=2
+  ad=750 pd=310 as=1500 ps=620
M1002 a_23_0# B a_7_0# w_n6_n6# pfet w=150 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 Y A gnd Gnd nfet w=20 l=2
+  ad=300 pd=150 as=300 ps=150
M1004 Y B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 Y C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a_7_0# a_23_0# 1.55fF
C1 A Y 0.05fF
C2 w_n6_n6# a_7_0# 0.32fF
C3 w_n6_n6# B 0.06fF
C4 a_23_0# Y 1.55fF
C5 C Y 0.24fF
C6 B a_7_0# 0.02fF
C7 w_n6_n6# Y 0.17fF
C8 w_n6_n6# vdd 0.17fF
C9 w_n6_n6# A 0.06fF
C10 Y gnd 1.21fF
C11 C a_23_0# 0.02fF
C12 A gnd 0.05fF
C13 vdd a_7_0# 1.55fF
C14 B Y 0.19fF
C15 w_n6_n6# a_23_0# 0.32fF
C16 w_n6_n6# C 0.06fF
C17 gnd Gnd 0.23fF
C18 Y Gnd 0.22fF
C19 a_23_0# Gnd 0.00fF
C20 a_7_0# Gnd 0.00fF
C21 vdd Gnd 0.01fF
C22 C Gnd 0.17fF
C23 B Gnd 0.17fF
C24 A Gnd 0.17fF
C25 w_n6_n6# Gnd 9.11fF
