magic
tech scmos
timestamp 1731236797
<< nwell >>
rect -6 -6 34 106
<< ntransistor >>
rect 5 -41 7 -21
rect 21 -41 23 -21
<< ptransistor >>
rect 5 0 7 100
rect 21 0 23 100
<< ndiffusion >>
rect 4 -41 5 -21
rect 7 -41 8 -21
rect 20 -41 21 -21
rect 23 -41 24 -21
<< pdiffusion >>
rect 4 0 5 100
rect 7 0 8 100
rect 20 0 21 100
rect 23 0 24 100
<< ndcontact >>
rect 0 -41 4 -21
rect 8 -41 12 -21
rect 16 -41 20 -21
rect 24 -41 28 -21
<< pdcontact >>
rect 0 0 4 100
rect 8 0 12 100
rect 16 0 20 100
rect 24 0 28 100
<< polysilicon >>
rect 5 100 7 103
rect 21 100 23 103
rect 5 -21 7 0
rect 21 -21 23 0
rect 5 -44 7 -41
rect 21 -44 23 -41
<< polycontact >>
rect 1 -18 5 -14
rect 17 -11 21 -7
<< metal1 >>
rect 0 100 4 109
rect 12 96 16 100
rect 13 -11 17 -7
rect 24 -14 28 0
rect -3 -18 1 -14
rect 8 -18 28 -14
rect 8 -21 12 -18
rect 24 -21 28 -18
rect 0 -46 4 -41
rect 16 -46 20 -41
rect 0 -50 20 -46
<< labels >>
rlabel metal1 10 -50 14 -46 1 gnd
rlabel metal1 24 -11 28 -7 1 Y
rlabel metal1 -3 -18 1 -14 1 A
rlabel metal1 13 -11 17 -7 1 B
rlabel metal1 0 105 4 109 5 vdd
<< end >>
