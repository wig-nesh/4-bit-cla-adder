magic
tech scmos
timestamp 1731231675
<< nwell >>
rect -6 -6 50 56
<< ntransistor >>
rect 5 -81 7 -21
rect 21 -81 23 -21
rect 37 -81 39 -21
<< ptransistor >>
rect 5 0 7 50
rect 21 0 23 50
rect 37 0 39 50
<< ndiffusion >>
rect 4 -81 5 -21
rect 7 -81 8 -21
rect 20 -81 21 -21
rect 23 -81 24 -21
rect 36 -81 37 -21
rect 39 -81 40 -21
<< pdiffusion >>
rect 4 0 5 50
rect 7 0 8 50
rect 20 0 21 50
rect 23 0 24 50
rect 36 0 37 50
rect 39 0 40 50
<< ndcontact >>
rect 0 -81 4 -21
rect 8 -81 12 -21
rect 16 -81 20 -21
rect 24 -81 28 -21
rect 32 -81 36 -21
rect 40 -81 44 -21
<< pdcontact >>
rect 0 0 4 50
rect 8 0 12 50
rect 16 0 20 50
rect 24 0 28 50
rect 32 0 36 50
rect 40 0 44 50
<< polysilicon >>
rect 5 50 7 53
rect 21 50 23 53
rect 37 50 39 53
rect 5 -21 7 0
rect 21 -21 23 0
rect 37 -21 39 0
rect 5 -84 7 -81
rect 21 -84 23 -81
rect 37 -84 39 -81
<< polycontact >>
rect 1 -11 5 -7
rect 17 -18 21 -14
rect 33 -18 37 -14
<< metal1 >>
rect 0 55 36 59
rect 0 50 4 55
rect 16 50 20 55
rect 32 50 36 55
rect 8 -7 12 0
rect 24 -7 28 0
rect 40 -7 44 0
rect -3 -11 1 -7
rect 8 -11 44 -7
rect 13 -18 17 -14
rect 29 -18 33 -14
rect 40 -21 44 -11
rect 12 -25 16 -21
rect 28 -25 32 -21
rect 0 -90 4 -81
<< labels >>
rlabel metal1 10 55 14 59 5 vdd
rlabel metal1 -3 -11 1 -7 1 A
rlabel metal1 13 -18 17 -14 1 B
rlabel metal1 29 -18 33 -14 1 C
rlabel metal1 40 -11 44 -7 1 Y
rlabel metal1 0 -90 4 -86 1 gnd
<< end >>
