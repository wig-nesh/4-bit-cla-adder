* .include ../../../tech_files/TSMC_180nm.txt

* .param SUPPLY=1.8
* .param LAMBDA=0.09u
* .param width_N={20*LAMBDA}
* .param width_P={2.5*width_N}
* .param length={2*LAMBDA}
* .global gnd vdd

* VDD vdd gnd SUPPLY
* vinA A gnd PULSE(0 SUPPLY 10ns 1ps 1ps 10ns 20ns)
* vinB B gnd PULSE(0 SUPPLY  5ns 1ps 1ps  5ns 10ns)

.subckt nor_cmos A B Y 
    .param width_P = 2*width_P
    MnA Y A gnd gnd CMOSN W={width_N} L={length} 
    + AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
    + AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
    MnB Y B gnd gnd CMOSN W={width_N} L={length} 
    + AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
    + AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
    MpA x A vdd vdd CMOSP W={width_P} L={length} 
    + AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} 
    + AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
    MpB Y B   x vdd CMOSP W={width_P} L={length} 
    + AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} 
    + AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
.ends

* Xand A B Y nor_cmos

* .tran 1n 20n 

* .measure tran t_in WHEN v(B)=0.5*SUPPLY CROSS=1
* .measure tran t_out WHEN v(Y)=0.5*SUPPLY CROSS=1
* .measure tran t_delay PARAM='t_out-t_in'

* .control
*     set hcopypscolor = 1
*     set color0=beige
*     set color1=black
*     set color2=blue
*     set color3=darkgreen
*     set color4=darkred
*     set color5=darkviolet
*     set color6=darkorange

*     run
*     plot v(A)+4 v(B)+2 v(Y)
* .endc