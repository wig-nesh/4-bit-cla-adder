magic
tech scmos
timestamp 1732120796
<< nwell >>
rect 997 318 1021 380
rect 997 98 1021 225
rect 997 -122 1021 4
<< ntransistor >>
rect 1008 290 1010 310
rect 1008 233 1010 253
rect 1008 70 1010 90
rect 1008 12 1010 32
rect 1008 -150 1010 -130
<< ptransistor >>
rect 1008 324 1010 374
rect 1008 169 1010 219
rect 1008 104 1010 154
rect 1008 -52 1010 -2
rect 1008 -116 1010 -66
<< ndiffusion >>
rect 1007 290 1008 310
rect 1010 290 1011 310
rect 1007 233 1008 253
rect 1010 233 1011 253
rect 1007 70 1008 90
rect 1010 70 1011 90
rect 1007 12 1008 32
rect 1010 12 1011 32
rect 1007 -150 1008 -130
rect 1010 -150 1011 -130
<< pdiffusion >>
rect 1007 324 1008 374
rect 1010 324 1011 374
rect 1007 169 1008 219
rect 1010 169 1011 219
rect 1007 104 1008 154
rect 1010 104 1011 154
rect 1007 -52 1008 -2
rect 1010 -52 1011 -2
rect 1007 -116 1008 -66
rect 1010 -116 1011 -66
<< ndcontact >>
rect 1003 290 1007 310
rect 1011 290 1015 310
rect 1003 233 1007 253
rect 1011 233 1015 253
rect 1003 70 1007 90
rect 1011 70 1015 90
rect 1003 12 1007 32
rect 1011 12 1015 32
rect 1003 -150 1007 -130
rect 1011 -150 1015 -130
<< pdcontact >>
rect 1003 324 1007 374
rect 1011 324 1015 374
rect 1003 169 1007 219
rect 1011 169 1015 219
rect 1003 104 1007 154
rect 1011 104 1015 154
rect 1003 -52 1007 -2
rect 1011 -52 1015 -2
rect 1003 -116 1007 -66
rect 1011 -116 1015 -66
<< polysilicon >>
rect 1008 374 1010 377
rect 1008 310 1010 324
rect 1008 287 1010 290
rect 1008 253 1010 256
rect 1008 219 1010 233
rect 1008 166 1010 169
rect 1008 154 1010 157
rect 1008 90 1010 104
rect 1008 67 1010 70
rect 1008 32 1010 35
rect 1008 -2 1010 12
rect 1008 -55 1010 -52
rect 1008 -66 1010 -63
rect 1008 -130 1010 -116
rect 1008 -153 1010 -150
<< polycontact >>
rect 1004 313 1008 317
rect 1004 226 1008 230
rect 1004 93 1008 97
rect 1004 5 1008 9
rect 1004 -127 1008 -123
<< metal1 >>
rect -179 408 52 412
rect -179 287 -175 408
rect 92 377 96 381
rect -106 335 19 339
rect -106 321 -102 335
rect 122 321 130 405
rect 156 377 160 381
rect 955 379 1007 383
rect 579 374 827 378
rect 955 377 959 379
rect 1003 374 1007 379
rect 579 367 583 374
rect 471 363 501 367
rect 553 363 579 367
rect 234 335 252 339
rect -38 315 18 319
rect 14 305 18 315
rect 14 302 20 305
rect -179 67 -175 285
rect 248 276 252 335
rect 248 272 267 276
rect 271 272 335 276
rect -74 253 -70 255
rect -148 243 -144 247
rect 248 231 252 272
rect 23 227 252 231
rect 331 256 335 272
rect 331 252 413 256
rect -172 209 -88 217
rect 51 203 55 227
rect 113 204 117 227
rect 175 205 179 227
rect 237 205 241 227
rect 331 209 335 252
rect 409 235 413 252
rect 471 235 475 363
rect 565 331 572 335
rect 1011 317 1015 324
rect 991 313 1004 317
rect 1011 313 1024 317
rect 923 307 926 311
rect 1011 310 1015 313
rect 1003 279 1007 290
rect 825 269 909 276
rect 959 275 1007 279
rect 583 267 909 269
rect 583 265 825 267
rect 409 231 475 235
rect -148 179 -144 183
rect -74 171 -70 174
rect 347 173 351 228
rect 409 209 413 231
rect 471 209 475 231
rect 425 173 429 187
rect 487 173 491 177
rect 67 169 71 173
rect 129 169 133 173
rect 191 169 195 173
rect 12 159 16 169
rect 74 159 78 169
rect 136 159 140 169
rect 198 160 202 170
rect 252 169 256 173
rect 260 115 264 173
rect 579 107 583 265
rect 1003 253 1007 275
rect 923 231 926 235
rect 1011 230 1015 233
rect 991 226 1004 230
rect 1011 226 1024 230
rect 1011 219 1015 226
rect 730 201 776 205
rect 780 201 815 205
rect 811 168 815 201
rect 754 162 765 166
rect 811 164 850 168
rect -72 103 53 107
rect 55 103 208 107
rect 241 103 727 107
rect -72 99 -38 103
rect 35 96 39 100
rect 97 96 101 100
rect 159 96 163 100
rect 221 96 225 100
rect -179 -77 -175 64
rect -74 32 -70 36
rect 33 33 35 35
rect 51 32 55 36
rect 113 32 117 36
rect 175 32 179 36
rect 237 32 241 36
rect 252 30 256 51
rect 261 33 265 37
rect -148 23 -144 27
rect 252 26 276 30
rect 363 13 367 37
rect 457 6 461 37
rect 535 9 539 37
rect 597 33 601 37
rect 23 0 209 4
rect -172 -11 -88 -3
rect 130 -36 134 0
rect -148 -41 -144 -37
rect -74 -49 -70 -47
rect 347 -62 351 1
rect 441 -42 445 2
rect 519 -21 523 1
rect 581 -21 585 1
rect 519 -25 549 -21
rect 553 -25 585 -21
rect 441 -44 471 -42
rect 519 -44 523 -25
rect 441 -46 499 -44
rect 441 -62 445 -46
rect 471 -48 499 -46
rect 526 -48 556 -44
rect 347 -66 445 -62
rect 6 -70 20 -66
rect -179 -173 -175 -81
rect 6 -109 10 -70
rect 84 -72 86 -68
rect 166 -72 168 -68
rect 347 -82 351 -66
rect 253 -86 351 -82
rect -38 -113 10 -109
rect -106 -125 -102 -114
rect -106 -129 19 -125
rect 92 -146 96 -142
rect 122 -170 130 -86
rect 253 -96 257 -86
rect 234 -100 257 -96
rect 315 -133 319 -86
rect 347 -107 351 -86
rect 552 -94 556 -48
rect 571 -98 600 -94
rect 347 -111 358 -107
rect 361 -111 464 -107
rect 389 -133 393 -111
rect 460 -133 464 -111
rect 156 -146 160 -142
rect -179 -176 52 -173
rect -179 -177 56 -176
rect 52 -250 56 -177
rect 124 -184 128 -170
rect 200 -177 204 -173
rect 228 -180 232 -170
rect 219 -184 232 -180
rect 596 -202 600 -98
rect 693 -97 697 103
rect 761 78 765 162
rect 925 163 959 165
rect 1003 163 1007 169
rect 925 159 1007 163
rect 925 157 959 159
rect 1003 154 1007 159
rect 1011 97 1015 104
rect 991 93 1004 97
rect 1011 93 1024 97
rect 923 87 926 91
rect 1011 90 1015 93
rect 761 74 767 78
rect 1003 59 1007 70
rect 959 55 1007 59
rect 825 46 909 55
rect 1003 32 1007 55
rect 923 11 926 15
rect 1011 9 1015 12
rect 991 5 1004 9
rect 1011 5 1024 9
rect 730 1 776 5
rect 779 1 811 5
rect 807 -52 811 1
rect 1011 -2 1015 5
rect 807 -56 843 -52
rect 925 -57 959 -55
rect 1003 -57 1007 -52
rect 925 -61 1007 -57
rect 925 -64 959 -61
rect 1003 -66 1007 -61
rect 693 -101 705 -97
rect 708 -101 769 -97
rect 1011 -123 1015 -116
rect 991 -127 1004 -123
rect 1011 -127 1024 -123
rect 923 -133 926 -129
rect 1011 -130 1015 -127
rect 690 -167 698 -163
rect 721 -179 725 -163
rect 751 -167 755 -153
rect 1003 -161 1007 -150
rect 781 -167 785 -163
rect 959 -165 1007 -161
rect 709 -197 766 -195
rect 705 -199 766 -197
rect 705 -202 709 -199
rect 596 -206 611 -202
rect 678 -206 709 -202
rect 113 -214 117 -210
rect 52 -254 83 -250
rect 267 -282 271 -234
rect 303 -235 460 -231
rect 464 -235 484 -231
rect 480 -249 484 -235
rect 480 -253 490 -249
rect 494 -253 552 -249
rect 223 -286 271 -282
<< m2contact >>
rect 83 302 88 307
rect 164 302 169 307
rect 11 154 16 159
rect 73 154 78 159
rect 135 154 140 159
rect 197 155 202 160
<< metal2 >>
rect 60 404 192 408
rect 195 404 826 408
rect 822 344 826 404
rect 347 331 494 335
rect 80 302 83 307
rect 169 302 172 307
rect -74 255 76 259
rect 72 178 76 255
rect 80 254 84 302
rect 168 254 172 302
rect 80 250 140 254
rect 168 250 202 254
rect 136 178 140 250
rect 198 178 202 250
rect 347 228 351 331
rect 425 323 511 327
rect 252 194 390 198
rect 0 174 35 178
rect 72 176 96 178
rect 136 176 158 178
rect 198 176 220 178
rect 72 174 97 176
rect 136 174 159 176
rect 198 174 221 176
rect 0 171 4 174
rect -74 167 4 171
rect 12 42 16 154
rect 31 96 35 174
rect 74 42 78 154
rect 93 96 97 174
rect 136 42 140 154
rect 155 96 159 174
rect 198 42 202 155
rect 217 96 221 174
rect 252 173 256 194
rect 260 186 358 190
rect 260 115 264 186
rect 252 111 264 115
rect 276 115 280 180
rect 292 124 296 180
rect 308 132 312 180
rect 354 170 358 186
rect 386 182 390 194
rect 425 187 429 323
rect 526 319 530 326
rect 487 315 530 319
rect 432 170 436 173
rect 354 166 436 170
rect 308 128 328 132
rect 292 120 312 124
rect 276 111 296 115
rect 252 54 256 111
rect 32 39 34 41
rect -74 35 11 39
rect 70 -11 74 33
rect 132 -11 136 32
rect 194 -11 198 32
rect 2 -15 74 -11
rect 80 -15 136 -11
rect 168 -15 198 -11
rect 2 -49 6 -15
rect -74 -53 6 -49
rect 80 -72 84 -15
rect 168 -72 172 -15
rect 292 -88 296 111
rect 260 -92 296 -88
rect 260 -165 264 -92
rect 308 -99 312 120
rect 276 -103 312 -99
rect 276 -162 280 -103
rect 324 -108 328 128
rect 386 21 390 166
rect 448 104 452 183
rect 487 177 491 315
rect 822 205 826 337
rect 765 147 769 164
rect 542 143 769 147
rect 448 100 500 104
rect 480 21 484 30
rect 386 17 484 21
rect 292 -112 328 -108
rect 61 -173 192 -169
rect 292 -186 296 -112
rect 363 -150 367 13
rect 496 -71 500 100
rect 542 36 546 143
rect 694 109 758 113
rect 597 33 656 37
rect 535 5 544 9
rect 496 -75 519 -71
rect 515 -87 519 -75
rect 540 -142 544 5
rect 540 -146 640 -142
rect 363 -154 608 -150
rect 437 -186 441 -161
rect 604 -172 608 -154
rect 636 -165 640 -146
rect 652 -165 656 33
rect 694 -186 698 109
rect 748 -1 752 98
rect 748 -4 755 -1
rect 751 -153 755 -4
rect 822 -18 826 202
rect 822 -95 826 -22
rect 849 -175 853 -135
rect 725 -179 853 -175
rect 234 -190 698 -186
rect 234 -222 238 -190
rect 195 -226 238 -222
<< metal3 >>
rect 595 331 606 335
rect 542 215 546 327
rect 129 211 562 215
rect 129 173 133 211
rect 191 199 452 203
rect 191 173 195 199
rect 276 191 374 195
rect 276 180 280 191
rect 370 165 374 191
rect 448 184 452 199
rect 386 174 390 180
rect 386 170 420 174
rect 370 161 406 165
rect 51 62 374 66
rect 51 36 55 62
rect 113 51 256 55
rect 113 36 117 51
rect 175 43 249 47
rect 175 36 179 43
rect 237 13 241 32
rect 245 21 249 43
rect 261 37 265 62
rect 292 21 296 26
rect 245 17 296 21
rect 308 13 312 26
rect 237 9 312 13
rect 370 16 374 62
rect 402 30 406 161
rect 416 26 420 170
rect 464 16 468 35
rect 542 16 546 36
rect 558 29 562 211
rect 602 133 606 331
rect 806 305 849 309
rect 806 167 810 305
rect 602 129 810 133
rect 806 105 810 129
rect 724 101 777 105
rect 785 97 808 101
rect 370 12 546 16
rect 331 -80 483 -76
rect 538 -80 697 -76
rect 260 -175 264 -168
rect 331 -169 335 -80
rect 499 -98 503 -87
rect 405 -102 503 -98
rect 405 -169 409 -102
rect 584 -130 597 -126
rect 545 -165 549 -130
rect 476 -169 549 -165
rect 350 -175 354 -169
rect 260 -179 354 -175
rect 593 -181 597 -130
rect 693 -170 697 -80
rect 728 -170 732 -166
rect 785 -167 789 97
rect 808 81 853 85
rect 808 33 812 81
rect 693 -174 732 -170
rect 758 -181 762 -167
rect 593 -185 762 -181
<< metal4 >>
rect 292 164 296 183
rect 715 164 719 170
rect 292 160 719 164
rect 256 51 719 55
rect 292 40 703 44
rect 292 26 296 40
rect 699 29 703 40
rect 715 37 719 51
rect 765 29 769 36
rect 699 25 769 29
<< metal5 >>
rect 935 313 991 317
rect 760 233 849 237
rect 67 218 576 222
rect 67 171 71 218
rect 571 116 576 218
rect 571 111 672 116
rect 416 -70 420 26
rect 457 -62 461 6
rect 457 -66 624 -62
rect 366 -74 565 -70
rect 276 -180 280 -159
rect 366 -162 370 -74
rect 561 -137 565 -74
rect 620 -166 624 -66
rect 668 -165 672 111
rect 760 85 764 233
rect 935 226 991 230
rect 935 93 991 97
rect 756 82 764 85
rect 756 33 760 82
rect 767 74 853 78
rect 849 17 853 74
rect 935 5 991 9
rect 935 -127 991 -123
rect 421 -180 425 -167
rect 276 -184 425 -180
<< pad >>
rect 493 331 498 336
rect 593 330 598 335
rect 510 323 515 328
rect 526 323 531 328
rect 542 323 547 328
rect 932 312 937 317
rect 989 313 994 318
rect 848 304 853 309
rect -76 254 -71 259
rect 848 233 853 238
rect 347 226 352 231
rect 933 225 938 230
rect 989 225 994 230
rect 425 185 430 190
rect 30 174 36 180
rect 92 174 98 180
rect 154 174 160 180
rect 215 174 221 180
rect 276 179 281 184
rect 292 179 297 184
rect 308 179 313 184
rect 370 179 375 184
rect 386 179 391 184
rect 448 180 453 185
rect -76 169 -71 174
rect 66 168 71 173
rect 128 169 133 174
rect 190 169 195 174
rect 251 169 256 174
rect 354 173 359 178
rect 432 172 437 177
rect 486 173 491 178
rect 805 168 810 173
rect 259 111 264 116
rect 754 107 759 112
rect 723 100 728 105
rect 775 101 780 106
rect 805 105 810 110
rect 31 95 36 100
rect 93 95 98 100
rect 155 95 160 100
rect 217 95 222 100
rect 748 95 753 100
rect 804 95 809 100
rect 933 92 938 97
rect 989 93 994 98
rect 848 81 853 86
rect 765 74 770 79
rect 252 50 257 55
rect -76 34 -71 39
rect 50 32 55 37
rect 112 32 117 37
rect 174 32 179 37
rect 236 31 241 36
rect 261 33 266 38
rect 370 33 375 38
rect 464 32 469 37
rect 542 32 547 37
rect 596 32 601 37
rect 755 33 760 38
rect 807 33 812 38
rect 292 25 297 30
rect 308 25 313 30
rect 324 25 329 30
rect 386 26 391 31
rect 402 26 407 31
rect 417 25 422 30
rect 480 25 485 30
rect 496 26 501 31
rect 558 26 563 31
rect 362 10 367 15
rect 848 13 853 18
rect 457 4 462 9
rect 535 5 540 10
rect 933 5 938 10
rect 989 4 994 9
rect -76 -50 -71 -45
rect 81 -74 86 -69
rect 167 -74 172 -69
rect 480 -81 485 -76
rect 534 -81 539 -76
rect 499 -88 504 -83
rect 515 -87 520 -82
rect 545 -131 550 -126
rect 582 -131 587 -126
rect 933 -128 938 -123
rect 989 -127 994 -122
rect 561 -137 566 -132
rect 848 -136 853 -131
rect 750 -156 755 -151
rect 276 -163 281 -158
rect 292 -163 297 -158
rect 366 -162 371 -157
rect 437 -163 442 -158
rect 260 -169 265 -164
rect 330 -169 335 -164
rect 350 -170 355 -165
rect 404 -169 409 -164
rect 421 -170 426 -165
rect 475 -169 480 -164
rect 620 -167 625 -162
rect 636 -167 641 -162
rect 652 -167 657 -162
rect 668 -168 673 -163
rect 728 -168 733 -163
rect 758 -168 763 -163
rect 784 -167 789 -162
rect 604 -174 609 -169
rect 721 -180 726 -175
rect 197 -227 202 -222
use pg_gen_optimized_unrouted  pg_gen_optimized_unrouted_0 ../../../ckt_blocks/pg_gen/optimized/post_layout
timestamp 1732120796
transform 1 0 4 0 1 1
box -4 -1 251 230
use d_ff_optimized  d_ff_optimized_2 ../../../ckt_blocks/d_ff/optimized/post_layout
timestamp 1732120796
transform 0 1 20 1 0 -140
box -37 -4 111 106
use d_ff_optimized  d_ff_optimized_3
timestamp 1732120796
transform 0 -1 232 1 0 -140
box -37 -4 111 106
use d_ff_optimized  d_ff_optimized_8
timestamp 1732120796
transform 1 0 119 0 1 -286
box -37 -4 111 106
use d_ff_optimized  d_ff_optimized_7
timestamp 1732120796
transform 1 0 -142 0 1 -113
box -37 -4 111 106
use d_ff_optimized  d_ff_optimized_6
timestamp 1732120796
transform 1 0 -142 0 -1 99
box -37 -4 111 106
use d_ff_optimized  d_ff_optimized_0
timestamp 1732120796
transform 0 -1 232 -1 0 375
box -37 -4 111 106
use d_ff_optimized  d_ff_optimized_5
timestamp 1732120796
transform 0 1 20 -1 0 375
box -37 -4 111 106
use d_ff_optimized  d_ff_optimized_4
timestamp 1732120796
transform 1 0 -142 0 -1 319
box -37 -4 111 106
use d_ff_optimized  d_ff_optimized_1
timestamp 1732120796
transform 1 0 -142 0 1 107
box -37 -4 111 106
use cla_gen_cmos_unrouted  cla_gen_cmos_unrouted_0 ../../../ckt_blocks/cla_gen/cmos/post_layout
timestamp 1732120796
transform 1 0 261 0 1 -85
box -1 -168 522 452
use d_ff_optimized  d_ff_optimized_10
timestamp 1732120796
transform 1 0 855 0 -1 157
box -37 -4 111 106
use d_ff_optimized  d_ff_optimized_11
timestamp 1732120796
transform 1 0 855 0 1 165
box -37 -4 111 106
use d_ff_optimized  d_ff_optimized_12
timestamp 1732120796
transform 1 0 855 0 -1 377
box -37 -4 111 106
use d_ff_optimized  d_ff_optimized_9
timestamp 1732120796
transform 1 0 855 0 1 -55
box -37 -4 111 106
use d_ff_optimized  d_ff_optimized_13
timestamp 1732120796
transform 1 0 855 0 -1 -63
box -37 -4 111 106
use sum_gen_optimized_unrouted  sum_gen_optimized_unrouted_0 ../../../ckt_blocks/sum_gen/optimized/post_layout
timestamp 1732120796
transform 1 0 711 0 1 1
box -4 0 99 204
<< labels >>
rlabel metal1 -10 -113 -6 -109 1 vdd
rlabel metal1 -10 -129 -6 -125 1 gnd
rlabel metal1 156 -146 160 -142 1 B0
rlabel metal1 92 -146 96 -142 1 B1
rlabel metal1 156 377 160 381 1 A0
rlabel metal1 92 377 96 381 1 A1
rlabel metal1 -148 -41 -144 -37 1 B2
rlabel metal1 -148 23 -144 27 1 B3
rlabel metal1 -148 179 -144 183 1 A3
rlabel metal1 -148 243 -144 247 1 A2
rlabel metal1 -11 -177 -7 -173 1 clk
rlabel metal1 113 -214 117 -210 1 C0
rlabel metal1 923 307 926 311 1 Q3s
rlabel metal1 923 231 926 235 1 Q2s
rlabel metal1 923 87 926 91 1 Q1s
rlabel metal1 923 11 926 15 1 Q0s
rlabel metal1 923 -133 926 -129 1 Qco
rlabel metal1 1019 313 1024 317 7 S3out
rlabel metal1 1019 226 1024 230 7 S2out
rlabel metal1 1019 93 1024 97 7 S1out
rlabel metal1 1019 5 1024 9 7 S0out
rlabel metal1 1019 -127 1024 -123 7 Cout
<< end >>
