* SPICE3 file created from nand_cmos.ext - technology: scmos

.option scale=0.09u

M1000 Y A vdd w_n6_n6# pfet w=50 l=2
+  ad=500 pd=220 as=500 ps=220
M1001 Y B vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 a_7_n41# A gnd Gnd nfet w=20 l=2
+  ad=200 pd=100 as=100 ps=50
M1003 Y B a_7_n41# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
C0 Y gnd 0.03fF
C1 B a_7_n41# 0.16fF
C2 vdd Y 1.64fF
C3 w_n6_n6# Y 0.15fF
C4 A vdd 0.02fF
C5 w_n6_n6# A 0.06fF
C6 gnd a_7_n41# 0.27fF
C7 B gnd 0.05fF
C8 A Y 0.05fF
C9 w_n6_n6# B 0.06fF
C10 Y a_7_n41# 0.21fF
C11 B Y 0.31fF
C12 w_n6_n6# vdd 0.19fF
C13 A B 0.27fF
