.include ../../../../tech_files/TSMC_180nm.txt

.param SUPPLY=1.8
.global gnd vdd

VDD vdd gnd SUPPLY
vinA A gnd PULSE(0 SUPPLY   20ns 1ps 1ps   20ns  40ns)
vinB B gnd PULSE(0 SUPPLY   10ns 1ps 1ps   10ns  20ns)
vinC C gnd PULSE(0 SUPPLY    5ns 1ps 1ps    5ns  10ns)
vinD D gnd PULSE(0 SUPPLY  2.5ns 1ps 1ps  2.5ns   5ns)
vinE E gnd PULSE(0 SUPPLY 1.25ns 1ps 1ps 1.25ns 2.5ns)

.option scale=0.09u

M1000 a_7_0# A vdd w_n6_n6# CMOSP w=250 l=2
+  ad=2500 pd=1020 as=1250 ps=510
M1001 a_39_0# C a_23_0# w_n6_n6# CMOSP w=250 l=2
+  ad=2500 pd=1020 as=2500 ps=1020
M1002 a_23_0# B a_7_0# w_n6_n6# CMOSP w=250 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 Y D gnd Gnd CMOSN w=20 l=2
+  ad=500 pd=250 as=500 ps=250
M1004 Y E gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 Y A gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 Y E a_55_0# w_n6_n6# CMOSP w=250 l=2
+  ad=1250 pd=510 as=2500 ps=1020
M1007 Y B gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 a_55_0# D a_39_0# w_n6_n6# CMOSP w=250 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 Y C gnd Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a_55_0# Y 2.58fF
C1 A gnd 0.05fF
C2 E a_55_0# 0.02fF
C3 a_7_0# a_23_0# 2.58fF
C4 D Y 0.19fF
C5 A Y 0.05fF
C6 w_n6_n6# a_39_0# 0.52fF
C7 B a_7_0# 0.02fF
C8 w_n6_n6# vdd 0.27fF
C9 w_n6_n6# C 0.06fF
C10 a_23_0# a_39_0# 2.58fF
C11 C Y 0.19fF
C12 w_n6_n6# Y 0.27fF
C13 C a_23_0# 0.02fF
C14 w_n6_n6# a_23_0# 0.52fF
C15 w_n6_n6# E 0.06fF
C16 w_n6_n6# B 0.06fF
C17 Y gnd 2.21fF
C18 a_39_0# a_55_0# 2.58fF
C19 E Y 0.24fF
C20 D a_39_0# 0.02fF
C21 vdd a_7_0# 2.58fF
C22 B Y 0.19fF
C23 w_n6_n6# a_55_0# 0.52fF
C24 w_n6_n6# a_7_0# 0.52fF
C25 w_n6_n6# D 0.06fF
C26 w_n6_n6# A 0.06fF
C27 gnd Gnd 0.41fF
C28 Y Gnd 0.38fF
C29 vdd Gnd 0.01fF
C30 E Gnd 0.17fF
C31 D Gnd 0.17fF
C32 C Gnd 0.17fF
C33 B Gnd 0.17fF
C34 A Gnd 0.17fF
C35 w_n6_n6# Gnd 23.16fF


.tran 1n 40n 

.measure tran t_in WHEN v(E)=0.5*SUPPLY CROSS=1
.measure tran t_out WHEN v(Y)=0.5*SUPPLY CROSS=1
.measure tran t_in1 WHEN v(A)=0.5*SUPPLY CROSS=2
.measure tran t_out1 WHEN v(Y)=0.5*SUPPLY CROSS=2
.measure tran t_delay10 PARAM='t_out-t_in'
.measure tran t_delay01 PARAM='t_out1-t_in1'

.control
    set hcopypscolor = 1
    set color0=beige
    set color1=black
    set color2=blue
    set color3=darkgreen
    set color4=darkred
    set color5=darkviolet
    set color6=darkorange

    run
    plot v(Y) v(E)+2 v(D)+4 v(C)+6 v(B)+8 v(A)+10
    set curplottitle="2023102019"
    hardcopy nor_5_cmos_post_tran.eps v(Y) v(E)+2 v(D)+4 v(C)+6 v(B)+8 v(A)+10
.endc
