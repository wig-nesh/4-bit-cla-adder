.include ../../../../tech_files/TSMC_180nm.txt

.param SUPPLY=1.8
.global gnd vdd

VDD vdd gnd SUPPLY
vinD     D gnd PULSE(0 SUPPLY  12ns 1ps 1ps  8ns 32ns)
vinClk clk gnd PULSE(0 SUPPLY   5ns 1ps 1ps   5ns 10ns)


.option scale=0.09u


.subckt inv_cmos IN w_0_0# gnd vdd OUT
M1000 OUT IN vdd w_0_0# CMOSP w=50 l=2
+  ad=250 pd=110 as=250 ps=110
M1001 OUT IN gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=100 ps=50
C0 OUT IN 0.05fF
C1 w_0_0# vdd 0.07fF
C2 OUT w_0_0# 0.07fF
C3 w_0_0# IN 0.06fF
C4 OUT gnd 0.21fF
C5 gnd IN 0.05fF
C6 OUT vdd 0.52fF
C7 IN vdd 0.02fF
C8 gnd Gnd 0.06fF
C9 OUT Gnd 0.05fF
C10 vdd Gnd 0.00fF
C11 IN Gnd 0.13fF
C12 w_0_0# Gnd 1.49fF
.ends


* Top level circuit d_ff_optimized

Xinv_cmos_3 inv_cmos_3/IN inv_cmos_4/w_0_0# gnd vdd inv_cmos_4/IN inv_cmos
Xinv_cmos_4 inv_cmos_4/IN inv_cmos_4/w_0_0# gnd vdd Q inv_cmos
Xinv_cmos_0 clk inv_cmos_0/w_0_0# gnd vdd inv_cmos_0/OUT inv_cmos
Xinv_cmos_1 inv_cmos_1/IN inv_cmos_2/w_0_0# gnd vdd inv_cmos_2/IN inv_cmos
Xinv_cmos_2 inv_cmos_2/IN inv_cmos_2/w_0_0# gnd vdd inv_cmos_2/OUT inv_cmos
M1000 Q inv_cmos_0/OUT inv_cmos_3/IN Gnd CMOSN w=20 l=2
+  ad=460 pd=50 as=122 ps=50
M1001 inv_cmos_2/OUT clk inv_cmos_3/IN Gnd CMOSN w=20 l=2
+  ad=720 pd=100 as=0 ps=0
M1002 inv_cmos_1/IN clk inv_cmos_2/OUT Gnd CMOSN w=20 l=2
+  ad=240 pd=32 as=0 ps=0
M1003 inv_cmos_1/IN inv_cmos_0/OUT D Gnd CMOSN w=20 l=2
+  ad=0 pd=0 as=100 ps=50
C0 inv_cmos_4/w_0_0# vdd 0.13fF
C1 inv_cmos_1/IN inv_cmos_2/IN 0.00fF
C2 gnd inv_cmos_2/OUT 0.03fF
C3 clk vdd 0.21fF
C4 inv_cmos_3/IN inv_cmos_4/IN 0.00fF
C5 inv_cmos_2/IN vdd 0.55fF
C6 Q vdd 0.68fF
C7 inv_cmos_1/IN vdd 0.26fF
C8 gnd inv_cmos_4/w_0_0# 0.01fF
C9 inv_cmos_2/OUT inv_cmos_0/OUT 0.05fF
C10 gnd inv_cmos_2/IN 0.23fF
C11 Q gnd 0.13fF
C12 gnd inv_cmos_1/IN 0.54fF
C13 inv_cmos_2/w_0_0# inv_cmos_2/OUT 0.01fF
C14 gnd vdd 0.06fF
C15 clk inv_cmos_0/OUT 0.39fF
C16 D inv_cmos_0/OUT 0.20fF
C17 inv_cmos_3/IN inv_cmos_2/OUT 0.21fF
C18 inv_cmos_2/IN inv_cmos_0/OUT 0.06fF
C19 inv_cmos_1/IN inv_cmos_0/OUT 0.07fF
C20 inv_cmos_4/w_0_0# inv_cmos_4/IN 0.00fF
C21 inv_cmos_4/w_0_0# inv_cmos_3/IN 0.04fF
C22 clk inv_cmos_2/w_0_0# 0.27fF
C23 inv_cmos_0/w_0_0# clk 0.10fF
C24 vdd inv_cmos_0/OUT 0.35fF
C25 clk inv_cmos_3/IN 0.05fF
C26 inv_cmos_2/IN inv_cmos_2/w_0_0# -0.00fF
C27 inv_cmos_1/IN inv_cmos_2/w_0_0# 0.03fF
C28 inv_cmos_3/IN inv_cmos_2/IN 0.00fF
C29 Q inv_cmos_3/IN 0.21fF
C30 inv_cmos_3/IN inv_cmos_1/IN 0.57fF
C31 inv_cmos_2/w_0_0# vdd 0.13fF
C32 inv_cmos_0/w_0_0# vdd 0.02fF
C33 gnd inv_cmos_0/OUT 0.03fF
C34 vdd inv_cmos_4/IN 0.55fF
C35 inv_cmos_3/IN vdd 0.50fF
C36 clk inv_cmos_2/OUT 0.33fF
C37 gnd inv_cmos_4/IN 0.24fF
C38 gnd inv_cmos_3/IN 0.60fF
C39 inv_cmos_2/IN inv_cmos_2/OUT 0.12fF
C40 inv_cmos_1/IN inv_cmos_2/OUT 0.35fF
C41 inv_cmos_2/w_0_0# inv_cmos_0/OUT 0.01fF
C42 inv_cmos_2/OUT vdd 0.58fF
C43 inv_cmos_0/w_0_0# inv_cmos_0/OUT 0.09fF
C44 clk inv_cmos_2/IN 0.09fF
C45 inv_cmos_3/IN inv_cmos_0/OUT 0.00fF
C46 clk inv_cmos_1/IN 0.19fF
C47 inv_cmos_1/IN D 0.21fF
C48 inv_cmos_0/OUT Gnd 0.33fF
C49 inv_cmos_4/IN Gnd -0.04fF
C50 vdd Gnd 0.26fF
C51 D Gnd 0.01fF
C52 inv_cmos_2/OUT Gnd 0.21fF
C53 inv_cmos_2/IN Gnd 0.01fF
C54 inv_cmos_1/IN Gnd 0.84fF
C55 gnd Gnd 0.42fF
C56 clk Gnd 0.77fF
C57 Q Gnd -0.04fF
C58 inv_cmos_3/IN Gnd 0.11fF
.end


.tran 1n 160n 

.measure tran t_in WHEN v(clk)=0.5*SUPPLY CROSS=3
.measure tran t_out WHEN v(Q)=0.5*SUPPLY CROSS=1
.measure tran t_delay PARAM='t_out-t_in'

.control
    set hcopypscolor = 1
    set color0=beige
    set color1=black
    set color2=blue
    set color3=darkgreen
    set color4=darkred
    set color5=darkviolet
    set color6=darkorange

    run
    plot v(clk)+4 v(D)+2 v(Q)
.endc
