* SPICE3 file created from nor_5_cmos.ext - technology: scmos

.option scale=0.09u

M1000 a_7_0# A vdd w_n6_n6# pfet w=250 l=2
+  ad=2500 pd=1020 as=1250 ps=510
M1001 a_39_0# C a_23_0# w_n6_n6# pfet w=250 l=2
+  ad=2500 pd=1020 as=2500 ps=1020
M1002 a_23_0# B a_7_0# w_n6_n6# pfet w=250 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 Y D gnd Gnd nfet w=20 l=2
+  ad=500 pd=250 as=500 ps=250
M1004 Y E gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 Y A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 Y E a_55_0# w_n6_n6# pfet w=250 l=2
+  ad=1250 pd=510 as=2500 ps=1020
M1007 Y B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 a_55_0# D a_39_0# w_n6_n6# pfet w=250 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 Y C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a_55_0# Y 2.58fF
C1 A gnd 0.05fF
C2 E a_55_0# 0.02fF
C3 a_7_0# a_23_0# 2.58fF
C4 D Y 0.19fF
C5 A Y 0.05fF
C6 w_n6_n6# a_39_0# 0.52fF
C7 B a_7_0# 0.02fF
C8 w_n6_n6# vdd 0.27fF
C9 w_n6_n6# C 0.06fF
C10 a_23_0# a_39_0# 2.58fF
C11 C Y 0.19fF
C12 w_n6_n6# Y 0.27fF
C13 C a_23_0# 0.02fF
C14 w_n6_n6# a_23_0# 0.52fF
C15 w_n6_n6# E 0.06fF
C16 w_n6_n6# B 0.06fF
C17 Y gnd 2.21fF
C18 a_39_0# a_55_0# 2.58fF
C19 E Y 0.24fF
C20 D a_39_0# 0.02fF
C21 vdd a_7_0# 2.58fF
C22 B Y 0.19fF
C23 w_n6_n6# a_55_0# 0.52fF
C24 w_n6_n6# a_7_0# 0.52fF
C25 w_n6_n6# D 0.06fF
C26 w_n6_n6# A 0.06fF
C27 gnd Gnd 0.41fF
C28 Y Gnd 0.38fF
C29 vdd Gnd 0.01fF
C30 E Gnd 0.17fF
C31 D Gnd 0.17fF
C32 C Gnd 0.17fF
C33 B Gnd 0.17fF
C34 A Gnd 0.17fF
C35 w_n6_n6# Gnd 23.16fF
