* SPICE3 file created from nand_4_cmos.ext - technology: scmos

.option scale=0.09u

M1000 Y D a_39_n101# Gnd nfet w=80 l=2
+  ad=400 pd=170 as=800 ps=340
M1001 Y A vdd w_n6_n6# pfet w=50 l=2
+  ad=1000 pd=440 as=1000 ps=440
M1002 Y C vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 Y B vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_7_n101# A gnd Gnd nfet w=80 l=2
+  ad=800 pd=340 as=400 ps=170
M1005 a_39_n101# C a_23_n101# Gnd nfet w=80 l=2
+  ad=0 pd=0 as=800 ps=340
M1006 a_23_n101# B a_7_n101# Gnd nfet w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 Y D vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a_7_n101# a_23_n101# 0.82fF
C1 a_23_n101# C 0.10fF
C2 Y A 0.05fF
C3 Y vdd 3.78fF
C4 A w_n6_n6# 0.06fF
C5 w_n6_n6# vdd 0.34fF
C6 a_23_n101# a_39_n101# 0.82fF
C7 D a_39_n101# 0.10fF
C8 a_7_n101# B 0.10fF
C9 Y C 0.19fF
C10 Y D 0.24fF
C11 C w_n6_n6# 0.06fF
C12 Y a_39_n101# 0.82fF
C13 D w_n6_n6# 0.06fF
C14 A vdd 0.02fF
C15 Y B 0.19fF
C16 a_7_n101# gnd 0.82fF
C17 Y w_n6_n6# 0.29fF
C18 B w_n6_n6# 0.06fF
