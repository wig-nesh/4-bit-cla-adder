* .include ../../../tech_files/TSMC_180nm.txt

* .param SUPPLY=1.8
* .param LAMBDA=0.09u
* .param width_N={20*LAMBDA}
* .param width_P={2.5*width_N}
* .param length={2*LAMBDA}
* .global gnd vdd

* VDD vdd gnd SUPPLY
* vinA A gnd PULSE(0 SUPPLY 10ns 1ps 1ps 10ns 20ns)

.subckt inv_cmos IN OUT
    Mn OUT IN gnd gnd CMOSN W={width_N} L={2*LAMBDA} 
    + AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
    + AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
    Mp OUT IN vdd vdd CMOSP W={width_P} L={2*LAMBDA} 
    + AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} 
    + AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
.ends

* Xinv A Y inv_cmos

* .tran 1n 20n 

* .measure tran t_in WHEN v(A)=0.5*SUPPLY CROSS=1
* .measure tran t_out WHEN v(Y)=0.5*SUPPLY CROSS=1
* .measure tran t_delay PARAM='t_out-t_in'

* .control
*     set hcopypscolor = 1
*     set color0=beige
*     set color1=black
*     set color2=blue
*     set color3=darkgreen
*     set color4=darkred
*     set color5=darkviolet
*     set color6=darkorange

*     run
*     plot v(A)+2 v(Y)
* .endc