magic
tech scmos
timestamp 1731798549
<< ntransistor >>
rect 65 73 67 93
rect -1 48 1 68
rect -1 9 1 29
rect 57 9 59 29
<< ndiffusion >>
rect 64 73 65 93
rect 67 73 68 93
rect -2 48 -1 68
rect 1 48 2 68
rect -2 9 -1 29
rect 1 9 2 29
rect 56 9 57 29
rect 59 9 60 29
<< ndcontact >>
rect 60 73 64 93
rect 68 73 72 93
rect -6 48 -2 68
rect 2 48 6 68
rect -6 9 -2 29
rect 2 9 6 29
rect 52 9 56 29
rect 60 9 64 29
<< polysilicon >>
rect 65 93 67 96
rect -1 68 1 71
rect 65 57 67 73
rect -1 40 1 48
rect -1 29 1 36
rect 57 29 59 48
rect -1 6 1 9
rect 57 6 59 9
<< polycontact >>
rect 61 59 65 63
rect -5 41 -1 45
rect 53 41 57 45
rect -5 32 -1 36
<< metal1 >>
rect 76 102 88 104
rect -26 98 54 102
rect 76 100 100 102
rect -6 68 -2 72
rect -14 45 -10 59
rect 51 56 54 98
rect 88 98 100 100
rect 60 93 64 95
rect 68 70 72 73
rect 68 66 76 70
rect 91 66 92 70
rect 57 59 61 63
rect 92 60 96 64
rect 51 53 73 56
rect -22 38 -18 42
rect -14 41 -5 45
rect 2 44 17 48
rect 56 45 57 49
rect -37 32 -34 36
rect -14 36 -10 41
rect 13 37 17 44
rect -18 32 -10 36
rect -5 36 -1 37
rect 32 32 33 36
rect 48 32 55 36
rect 2 29 6 32
rect 52 29 56 32
rect -6 6 -2 9
rect 60 7 64 9
rect -30 2 40 3
rect 70 4 73 53
rect -30 -1 44 2
rect 70 0 84 4
rect 88 0 100 4
rect 36 -2 44 -1
<< m2contact >>
rect 59 95 64 100
rect 51 45 56 50
rect -34 32 -29 37
rect 13 32 18 37
rect 60 2 65 7
<< metal2 >>
rect 64 96 111 100
rect 107 68 111 96
rect 49 45 51 49
rect 5 41 53 45
rect -33 37 9 41
rect -9 32 -5 37
rect 13 6 17 32
rect 13 2 60 6
<< metal3 >>
rect -14 59 59 63
rect 2 37 56 40
rect 2 36 55 37
rect 2 32 6 36
rect 107 8 111 68
rect -6 4 111 8
<< metal5 >>
rect 72 2 76 104
rect 44 -2 76 2
<< pad >>
rect 72 101 77 106
rect 106 67 111 72
rect -14 58 -9 63
rect 56 58 61 63
rect -9 32 -4 37
rect 2 31 7 36
rect 51 32 56 37
rect -7 4 -2 9
rect 42 -4 47 1
use inv_cmos  inv_cmos_0 ../../../inv/cmos/post_layout
timestamp 1731226851
transform 1 0 -36 0 1 37
box 0 -37 24 65
use inv_cmos  inv_cmos_1
timestamp 1731226851
transform 1 0 14 0 1 37
box 0 -37 24 65
use inv_cmos  inv_cmos_2
timestamp 1731226851
transform 1 0 30 0 1 37
box 0 -37 24 65
use inv_cmos  inv_cmos_4
timestamp 1731226851
transform -1 0 94 0 -1 65
box 0 -37 24 65
use inv_cmos  inv_cmos_3
timestamp 1731226851
transform -1 0 110 0 -1 65
box 0 -37 24 65
<< labels >>
rlabel metal1 -37 32 -33 36 3 clk
rlabel metal1 -6 68 -2 72 1 D
rlabel metal1 -7 98 -3 102 1 vdd
rlabel metal1 -15 -1 -11 3 1 gnd
rlabel metal1 68 66 71 70 1 Q
<< end >>
