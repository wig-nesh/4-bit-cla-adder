.include ../../../../tech_files/TSMC_180nm.txt

.param SUPPLY=1.8
.global gnd vdd

VDD vdd gnd SUPPLY
vinA A gnd PULSE(0 SUPPLY 10ns 1ps 1ps 10ns 20ns)
vinB B gnd PULSE(0 SUPPLY  5ns 1ps 1ps  5ns 10ns)

.option scale=0.09u

M1000 Y A vdd w_n6_n6# CMOSP w=50 l=2
+  ad=500 pd=220 as=500 ps=220
M1001 Y B vdd w_n6_n6# CMOSP w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 a_7_n41# A gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=100 ps=50
M1003 Y B a_7_n41# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
C0 Y gnd 0.03fF
C1 B a_7_n41# 0.16fF
C2 vdd Y 1.64fF
C3 w_n6_n6# Y 0.15fF
C4 A vdd 0.02fF
C5 w_n6_n6# A 0.06fF
C6 gnd a_7_n41# 0.27fF
C7 B gnd 0.05fF
C8 A Y 0.05fF
C9 w_n6_n6# B 0.06fF
C10 Y a_7_n41# 0.21fF
C11 B Y 0.31fF
C12 w_n6_n6# vdd 0.19fF
C13 A B 0.27fF



.tran 1n 20n 

.measure tran t_in WHEN v(B)=0.5*SUPPLY CROSS=3
.measure tran t_out WHEN v(Y)=0.5*SUPPLY CROSS=1
.measure tran t_delay PARAM='t_out-t_in'

.control
    set hcopypscolor = 1
    set color0=beige
    set color1=black
    set color2=blue
    set color3=darkgreen
    set color4=darkred
    set color5=darkviolet
    set color6=darkorange

    run
    plot v(A)+4 v(B)+2 v(Y)
.endc