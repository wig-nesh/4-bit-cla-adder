* SPICE3 file created from nor_4_cmos.ext - technology: scmos

.option scale=0.09u

M1000 Y D gnd Gnd nfet w=20 l=2
+  ad=400 pd=200 as=400 ps=200
M1001 a_7_0# A vdd w_n6_n6# pfet w=200 l=2
+  ad=2000 pd=820 as=1000 ps=410
M1002 a_39_0# C a_23_0# w_n6_n6# pfet w=200 l=2
+  ad=2000 pd=820 as=2000 ps=820
M1003 a_23_0# B a_7_0# w_n6_n6# pfet w=200 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 Y A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 Y B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 Y C gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 Y D a_39_0# w_n6_n6# pfet w=200 l=2
+  ad=1000 pd=410 as=0 ps=0
C0 a_23_0# a_39_0# 2.06fF
C1 C Y 0.19fF
C2 w_n6_n6# Y 0.22fF
C3 w_n6_n6# a_7_0# 0.42fF
C4 w_n6_n6# C 0.06fF
C5 a_39_0# Y 2.06fF
C6 A gnd 0.05fF
C7 vdd a_7_0# 2.06fF
C8 B Y 0.19fF
C9 w_n6_n6# a_39_0# 0.42fF
C10 w_n6_n6# vdd 0.22fF
C11 w_n6_n6# B 0.06fF
C12 Y gnd 1.71fF
C13 a_7_0# a_23_0# 2.06fF
C14 D Y 0.24fF
C15 A Y 0.05fF
C16 w_n6_n6# a_23_0# 0.42fF
C17 w_n6_n6# D 0.06fF
C18 w_n6_n6# A 0.06fF
C19 gnd Gnd 0.32fF
C20 Y Gnd 0.30fF
C21 a_39_0# Gnd 0.00fF
C22 a_23_0# Gnd 0.00fF
C23 a_7_0# Gnd 0.00fF
C24 vdd Gnd 0.01fF
C25 D Gnd 0.17fF
C26 C Gnd 0.17fF
C27 B Gnd 0.17fF
C28 A Gnd 0.17fF
C29 w_n6_n6# Gnd 15.33fF
