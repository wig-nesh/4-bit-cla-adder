.include ../../../../tech_files/TSMC_180nm.txt

.param SUPPLY=1.8
.param LAMBDA=0.09u
.global gnd vdd

VDD vdd gnd SUPPLY
vinA A gnd PULSE(0 SUPPLY   20ns 1ps 1ps   20ns  40ns)
vinB B gnd PULSE(0 SUPPLY   10ns 1ps 1ps   10ns  20ns)
vinC C gnd PULSE(0 SUPPLY    5ns 1ps 1ps    5ns  10ns)
vinD D gnd PULSE(0 SUPPLY  2.5ns 1ps 1ps  2.5ns   5ns)
vinE E gnd PULSE(0 SUPPLY 1.25ns 1ps 1ps 1.25ns 2.5ns)

.option scale=0.09u

M1000 Y A vdd w_n6_n6# CMOSP w=50 l=2
+  ad=1250 pd=550 as=1250 ps=550
M1001 Y C vdd w_n6_n6# CMOSP w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 Y B vdd w_n6_n6# CMOSP w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 Y E a_55_n121# Gnd CMOSN w=100 l=2
+  ad=500 pd=210 as=1000 ps=420
M1004 a_55_n121# D a_39_n121# Gnd CMOSN w=100 l=2
+  ad=0 pd=0 as=1000 ps=420
M1005 Y E vdd w_n6_n6# CMOSP w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 Y D vdd w_n6_n6# CMOSP w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_7_n121# A gnd Gnd CMOSN w=100 l=2
+  ad=1000 pd=420 as=500 ps=210
M1008 a_39_n121# C a_23_n121# Gnd CMOSN w=100 l=2
+  ad=0 pd=0 as=1000 ps=420
M1009 a_23_n121# B a_7_n121# Gnd CMOSN w=100 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_n6_n6# C 0.06fF
C1 gnd a_7_n121# 1.03fF
C2 B a_7_n121# 0.10fF
C3 D Y 0.19fF
C4 A Y 0.05fF
C5 a_39_n121# a_55_n121# 1.03fF
C6 w_n6_n6# E 0.06fF
C7 w_n6_n6# B 0.06fF
C8 E a_55_n121# 0.10fF
C9 a_7_n121# a_23_n121# 1.03fF
C10 C a_23_n121# 0.10fF
C11 vdd Y 4.87fF
C12 C Y 0.19fF
C13 w_n6_n6# Y 0.37fF
C14 A vdd 0.02fF
C15 w_n6_n6# D 0.06fF
C16 Y a_55_n121# 1.03fF
C17 w_n6_n6# A 0.06fF
C18 a_23_n121# a_39_n121# 1.03fF
C19 D a_39_n121# 0.10fF
C20 E Y 0.24fF
C21 B Y 0.19fF
C22 w_n6_n6# vdd 0.42fF


Xnand A B C D E Y nand_5_cmos

.tran 1n 40n 

.measure tran t_in WHEN v(E)=0.5*SUPPLY CROSS=31
.measure tran t_out WHEN v(Y)=0.5*SUPPLY CROSS=1
.measure tran t_delay PARAM='t_out-t_in'

.control
    set hcopypscolor = 1
    set color0=beige
    set color1=black
    set color2=blue
    set color3=darkgreen
    set color4=darkred
    set color5=darkviolet
    set color6=darkorange

    run
    plot v(Y) v(E)+2 v(D)+4 v(C)+6 v(B)+8 v(A)+10
.endc
