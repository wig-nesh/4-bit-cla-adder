magic
tech scmos
timestamp 1731239310
<< nwell >>
rect -6 -6 66 56
<< ntransistor >>
rect 5 -101 7 -21
rect 21 -101 23 -21
rect 37 -101 39 -21
rect 53 -101 55 -21
<< ptransistor >>
rect 5 0 7 50
rect 21 0 23 50
rect 37 0 39 50
rect 53 0 55 50
<< ndiffusion >>
rect 4 -101 5 -21
rect 7 -101 8 -21
rect 20 -101 21 -21
rect 23 -101 24 -21
rect 36 -101 37 -21
rect 39 -101 40 -21
rect 52 -101 53 -21
rect 55 -101 56 -21
<< pdiffusion >>
rect 4 0 5 50
rect 7 0 8 50
rect 20 0 21 50
rect 23 0 24 50
rect 36 0 37 50
rect 39 0 40 50
rect 52 0 53 50
rect 55 0 56 50
<< ndcontact >>
rect 0 -101 4 -21
rect 8 -101 12 -21
rect 16 -101 20 -21
rect 24 -101 28 -21
rect 32 -101 36 -21
rect 40 -101 44 -21
rect 48 -101 52 -21
rect 56 -101 60 -21
<< pdcontact >>
rect 0 0 4 50
rect 8 0 12 50
rect 16 0 20 50
rect 24 0 28 50
rect 32 0 36 50
rect 40 0 44 50
rect 48 0 52 50
rect 56 0 60 50
<< polysilicon >>
rect 5 50 7 53
rect 21 50 23 53
rect 37 50 39 53
rect 53 50 55 53
rect 5 -21 7 0
rect 21 -21 23 0
rect 37 -21 39 0
rect 53 -21 55 0
rect 5 -104 7 -101
rect 21 -104 23 -101
rect 37 -104 39 -101
rect 53 -104 55 -101
<< polycontact >>
rect 1 -11 5 -7
rect 17 -18 21 -14
rect 33 -18 37 -14
rect 49 -18 53 -14
<< metal1 >>
rect 0 55 52 59
rect 0 50 4 55
rect 16 50 20 55
rect 32 50 36 55
rect 48 50 52 55
rect 8 -7 12 0
rect 24 -7 28 0
rect 40 -7 44 0
rect 56 -7 60 0
rect -3 -11 1 -7
rect 8 -11 60 -7
rect 13 -18 17 -14
rect 29 -18 33 -14
rect 45 -18 49 -14
rect 56 -21 60 -11
rect 12 -25 16 -21
rect 28 -25 32 -21
rect 44 -25 48 -21
rect 0 -110 4 -101
<< labels >>
rlabel metal1 10 55 14 59 5 vdd
rlabel metal1 -3 -11 1 -7 1 A
rlabel metal1 13 -18 17 -14 1 B
rlabel metal1 29 -18 33 -14 1 C
rlabel metal1 45 -18 49 -14 1 D
rlabel metal1 0 -110 4 -106 1 gnd
<< end >>
