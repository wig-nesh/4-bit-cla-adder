magic
tech scmos
timestamp 1731238409
<< nwell >>
rect -6 -6 34 56
<< ntransistor >>
rect 5 -61 7 -21
rect 21 -61 23 -21
<< ptransistor >>
rect 5 0 7 50
rect 21 0 23 50
<< ndiffusion >>
rect 4 -61 5 -21
rect 7 -61 8 -21
rect 20 -61 21 -21
rect 23 -61 24 -21
<< pdiffusion >>
rect 4 0 5 50
rect 7 0 8 50
rect 20 0 21 50
rect 23 0 24 50
<< ndcontact >>
rect 0 -61 4 -21
rect 8 -61 12 -21
rect 16 -61 20 -21
rect 24 -61 28 -21
<< pdcontact >>
rect 0 0 4 50
rect 8 0 12 50
rect 16 0 20 50
rect 24 0 28 50
<< polysilicon >>
rect 5 50 7 53
rect 21 50 23 53
rect 5 -21 7 0
rect 21 -21 23 0
rect 5 -64 7 -61
rect 21 -64 23 -61
<< polycontact >>
rect 1 -11 5 -7
rect 17 -18 21 -14
<< metal1 >>
rect 0 55 20 59
rect 0 50 4 55
rect 16 50 20 55
rect 8 -7 12 0
rect 24 -7 28 0
rect -3 -11 1 -7
rect 8 -11 28 -7
rect 13 -18 17 -14
rect 24 -21 28 -11
rect 0 -69 4 -61
rect 8 -65 20 -61
<< labels >>
rlabel metal1 10 55 14 59 5 vdd
rlabel metal1 24 -11 28 -7 1 Y
rlabel metal1 -3 -11 1 -7 1 A
rlabel metal1 13 -18 17 -14 1 B
rlabel metal1 0 -69 4 -65 1 gnd
<< end >>
