* .include ../../../tech_files/TSMC_180nm.txt
.include ../../inv/cmos/inv_cmos.cir

* .param SUPPLY=1.8
* .param LAMBDA=0.09u
* .param width_N={20*LAMBDA}
* .param width_P={2.5*width_N}
* .param length={2*LAMBDA}
* .global gnd vdd

* VDD vdd gnd SUPPLY
* vinD     D gnd PULSE(0 SUPPLY  12ns 1ps 1ps  8ns 32ns)
* vinClk clk gnd PULSE(0 SUPPLY   5ns 1ps 1ps   5ns 10ns)

.subckt d_ff_optimized D clk Q x z a
    Xinv1 clk clki inv_cmos
    Mn1 D clki x gnd CMOSN W={width_N} L={2*LAMBDA} 
    + AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
    + AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
    Xinv2 x z inv_cmos
    Xinv3 z y inv_cmos
    Mn2 x clk y gnd CMOSN W={width_N} L={2*LAMBDA} 
    + AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
    + AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
    Mn3 z clk a gnd CMOSN W={width_N} L={2*LAMBDA} 
    + AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
    + AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
    Mn4 a clki b gnd CMOSN W={width_N} L={2*LAMBDA} 
    + AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
    + AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
    Xinv4 a Q inv_cmos
    Xinv5 Q b inv_cmos
.ends


* Xdff D clk Q x z a d_ff_optimized

* .tran 1n 160n 

* .measure tran t_clk WHEN v(clk)=0.5*SUPPLY CROSS=3
* .measure tran t_q WHEN v(Q)=0.5*SUPPLY CROSS=1

* .measure tran t_m1_rise_l WHEN v(x)=0.1*1.2 CROSS=3
* .measure tran t_m1_rise_h WHEN v(x)=0.9*1.2 CROSS=1
* .measure tran t_m1_prop WHEN v(x)=0.5*1.2 CROSS=1
* .measure tran t_inv1_prop WHEN v(z)=0.5*SUPPLY CROSS=1

* .measure tran t_m2_fall_l WHEN v(z)=0.1*SUPPLY CROSS=1
* .measure tran t_m2_fall_h WHEN v(z)=0.9*SUPPLY CROSS=1
* .measure tran t_m2_prop WHEN v(a)=0.5*SUPPLY CROSS=1
* .measure tran t_inv2_prop WHEN v(Q)=0.5*SUPPLY CROSS=1

* .measure tran t_cq PARAM='t_q-t_clk'
* .measure tran t_su PARAM='t_m1_rise_h-t_m1_rise_l+t_inv1_prop-t_m1_prop'
* .measure tran t_h PARAM='t_m2_fall_l-t_m2_fall_h+t_inv2_prop-t_m2_prop'

* .control
*     set hcopypscolor = 1
*     set color0=beige
*     set color1=black
*     set color2=blue
*     set color3=darkgreen
*     set color4=darkred
*     set color5=darkviolet
*     set color6=darkorange

*     run
*     plot v(clk)+4 v(D)+2 v(Q)
*     set curplottitle="2023102019"
*     hardcopy d_ff_optimized_tran.eps v(clk)+4 v(D)+2 v(Q)
* .endc