* SPICE3 file created from xor_optimized.ext - technology: scmos

.option scale=0.09u

.global Vdd Gnd 

.subckt inv_cmos IN w_0_0# OUT
M1000 OUT IN vdd w_0_0# pfet w=50 l=2
+  ad=250 pd=110 as=250 ps=110
M1001 OUT IN gnd Gnd nfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
C0 IN vdd 0.02fF
C1 vdd w_0_0# 0.07fF
C2 OUT gnd 0.21fF
C3 IN gnd 0.05fF
C4 OUT IN 0.05fF
C5 OUT w_0_0# 0.07fF
C6 IN w_0_0# 0.06fF
C7 OUT vdd 0.52fF
C8 gnd Gnd 0.06fF
C9 OUT Gnd 0.05fF
C10 vdd Gnd 0.00fF
C11 IN Gnd 0.13fF
C12 w_0_0# Gnd 1.49fF
.ends


* Top level circuit xor_optimized

Xinv_cmos_0 B w_26_37# inv_cmos_0/OUT inv_cmos
M1000 Y A inv_cmos_0/OUT Gnd nfet w=20 l=2
+  ad=100 pd=50 as=100 ps=50
M1001 Y A B w_26_37# pfet w=50 l=2
+  ad=250 pd=110 as=320 ps=110
C0 w_26_37# Y 0.07fF
C1 A B 0.05fF
C2 inv_cmos_0/OUT B 0.70fF
C3 A w_26_37# 0.10fF
C4 inv_cmos_0/OUT Y 0.28fF
C5 B w_26_37# 0.28fF
C6 B Y 0.56fF
C7 Y Gnd 0.05fF
C8 A Gnd 0.01fF
C9 inv_cmos_0/OUT Gnd 0.06fF
C10 B Gnd 0.32fF
C11 w_26_37# Gnd 1.12fF
.end

