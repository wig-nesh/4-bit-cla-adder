.include ../../../tech_files/TSMC_180nm.txt

.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={20*LAMBDA}
.param width_P={2.5*width_N}
.param length={2*LAMBDA}
.global gnd vdd

VDD vdd gnd SUPPLY
vinD     D gnd PULSE(0 SUPPLY  12ns 1ps 1ps  8ns 32ns)
vinClk clk gnd PULSE(0 SUPPLY   5ns 1ps 1ps   5ns 10ns)

.subckt d_ff_cmos D clk Q Qi
    .subckt inv_cmos IN OUT
        Mn OUT IN gnd gnd CMOSN W={width_N} L={2*LAMBDA} 
        + AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
        + AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
        Mp OUT IN vdd vdd CMOSP W={width_P} L={2*LAMBDA} 
        + AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} 
        + AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
    .ends INV
    .subckt nand_cmos A B Y 
        MnA Y A   x gnd CMOSN W={width_N} L={length} 
        + AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
        + AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
        MnB x B gnd gnd CMOSN W={width_N} L={length} 
        + AS={5*width_N*LAMBDA} PS={10*LAMBDA+2*width_N} 
        + AD={5*width_N*LAMBDA} PD={10*LAMBDA+2*width_N}
        MpA Y A vdd vdd CMOSP W={width_P} L={length} 
        + AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} 
        + AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
        MpB Y B vdd vdd CMOSP W={width_P} L={length} 
        + AS={5*width_P*LAMBDA} PS={10*LAMBDA+2*width_P} 
        + AD={5*width_P*LAMBDA} PD={10*LAMBDA+2*width_P}
    .ends
    Xinv    D     Di inv_cmos
    Xnand1  D clk  x nand_cmos
    Xnand2 Di clk  y nand_cmos
    Xnand3  x  Qi  Q nand_cmos
    Xnand4  y   Q Qi nand_cmos
.ends

Xdff D clk Q Qi d_ff_cmos

.tran 1n 80n 

.measure tran t_in WHEN v(clk)=0.5*SUPPLY CROSS=3
.measure tran t_out WHEN v(Q)=0.5*SUPPLY CROSS=2
.measure tran t_delay PARAM='t_out-t_in'

.control
    set hcopypscolor = 1
    set color0=beige
    set color1=black
    set color2=blue
    set color3=darkgreen
    set color4=darkred
    set color5=darkviolet
    set color6=darkorange

    run
    plot v(clk)+4 v(D)+2 v(Q) V(Qi)-2
.endc