magic
tech scmos
timestamp 1731232449
<< nwell >>
rect -6 -6 82 56
<< ntransistor >>
rect 5 -121 7 -21
rect 21 -121 23 -21
rect 37 -121 39 -21
rect 53 -121 55 -21
rect 69 -121 71 -21
<< ptransistor >>
rect 5 0 7 50
rect 21 0 23 50
rect 37 0 39 50
rect 53 0 55 50
rect 69 0 71 50
<< ndiffusion >>
rect 4 -121 5 -21
rect 7 -121 8 -21
rect 20 -121 21 -21
rect 23 -121 24 -21
rect 36 -121 37 -21
rect 39 -121 40 -21
rect 52 -121 53 -21
rect 55 -121 56 -21
rect 68 -121 69 -21
rect 71 -121 72 -21
<< pdiffusion >>
rect 4 0 5 50
rect 7 0 8 50
rect 20 0 21 50
rect 23 0 24 50
rect 36 0 37 50
rect 39 0 40 50
rect 52 0 53 50
rect 55 0 56 50
rect 68 0 69 50
rect 71 0 72 50
<< ndcontact >>
rect 0 -121 4 -21
rect 8 -121 12 -21
rect 16 -121 20 -21
rect 24 -121 28 -21
rect 32 -121 36 -21
rect 40 -121 44 -21
rect 48 -121 52 -21
rect 56 -121 60 -21
rect 64 -121 68 -21
rect 72 -121 76 -21
<< pdcontact >>
rect 0 0 4 50
rect 8 0 12 50
rect 16 0 20 50
rect 24 0 28 50
rect 32 0 36 50
rect 40 0 44 50
rect 48 0 52 50
rect 56 0 60 50
rect 64 0 68 50
rect 72 0 76 50
<< polysilicon >>
rect 5 50 7 53
rect 21 50 23 53
rect 37 50 39 53
rect 53 50 55 53
rect 69 50 71 53
rect 5 -21 7 0
rect 21 -21 23 0
rect 37 -21 39 0
rect 53 -21 55 0
rect 69 -21 71 0
rect 5 -124 7 -121
rect 21 -124 23 -121
rect 37 -124 39 -121
rect 53 -124 55 -121
rect 69 -124 71 -121
<< polycontact >>
rect 1 -11 5 -7
rect 17 -18 21 -14
rect 33 -18 37 -14
rect 49 -18 53 -14
rect 65 -18 69 -14
<< metal1 >>
rect 0 55 68 59
rect 0 50 4 55
rect 16 50 20 55
rect 32 50 36 55
rect 48 50 52 55
rect 64 50 68 55
rect 8 -7 12 0
rect 24 -7 28 0
rect 40 -7 44 0
rect 56 -7 60 0
rect 72 -7 76 0
rect -3 -11 1 -7
rect 8 -11 76 -7
rect 13 -18 17 -14
rect 29 -18 33 -14
rect 45 -18 49 -14
rect 61 -18 65 -14
rect 72 -21 76 -11
rect 12 -25 16 -21
rect 28 -25 32 -21
rect 44 -25 48 -21
rect 60 -25 64 -21
rect 0 -130 4 -121
<< labels >>
rlabel metal1 10 55 14 59 5 vdd
rlabel metal1 -3 -11 1 -7 1 A
rlabel metal1 61 -18 65 -14 1 E
rlabel metal1 45 -18 49 -14 1 D
rlabel metal1 13 -18 17 -14 1 B
rlabel metal1 29 -18 33 -14 1 C
rlabel metal1 72 -11 76 -7 1 Y
rlabel metal1 0 -130 4 -126 1 gnd
<< end >>
