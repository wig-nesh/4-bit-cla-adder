* SPICE3 file created from nand_4_cmos.ext - technology: scmos

.option scale=0.09u

M1000 a_7_0# D a_39_n101# Gnd nfet w=80 l=2
+  ad=400 pd=170 as=800 ps=340
M1001 a_7_0# A vdd w_n6_n6# pfet w=50 l=2
+  ad=1000 pd=440 as=1000 ps=440
M1002 a_7_0# C vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_7_0# B vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_7_n101# A gnd Gnd nfet w=80 l=2
+  ad=800 pd=340 as=400 ps=170
M1005 a_39_n101# C a_23_n101# Gnd nfet w=80 l=2
+  ad=0 pd=0 as=800 ps=340
M1006 a_23_n101# B a_7_n101# Gnd nfet w=80 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 a_7_0# D vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a_7_0# a_39_n101# 0.82fF
C1 a_23_n101# C 0.10fF
C2 D a_39_n101# 0.10fF
C3 a_7_0# vdd 3.78fF
C4 a_7_0# A 0.05fF
C5 C w_n6_n6# 0.06fF
C6 B w_n6_n6# 0.06fF
C7 a_7_0# w_n6_n6# 0.29fF
C8 a_7_n101# gnd 0.82fF
C9 D w_n6_n6# 0.06fF
C10 a_23_n101# a_7_n101# 0.82fF
C11 a_7_0# C 0.19fF
C12 a_23_n101# a_39_n101# 0.82fF
C13 a_7_0# B 0.19fF
C14 D a_7_0# 0.24fF
C15 vdd A 0.02fF
C16 a_7_n101# B 0.10fF
C17 vdd w_n6_n6# 0.34fF
C18 A w_n6_n6# 0.06fF
