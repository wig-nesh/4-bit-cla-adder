.include ../../../../tech_files/TSMC_180nm.txt

.param SUPPLY=1.8
.global gnd vdd

VDD vdd gnd SUPPLY
vinA A gnd PULSE(0 SUPPLY 10ns 1ps 1ps 10ns 20ns)
vinB B gnd PULSE(0 SUPPLY  5ns 1ps 1ps  5ns 10ns)

.option scale=0.09u

M1000 a_7_n61# A gnd Gnd CMOSN w=40 l=2
+  ad=400 pd=180 as=200 ps=90
M1001 Y B a_7_n61# Gnd CMOSN w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1002 Y A vdd w_n6_n6# CMOSP w=50 l=2
+  ad=500 pd=220 as=500 ps=220
M1003 Y B vdd w_n6_n6# CMOSP w=50 l=2
+  ad=0 pd=0 as=0 ps=0
C0 a_7_n61# Y 0.41fF
C1 A vdd 0.02fF
C2 w_n6_n6# vdd 0.16fF
C3 A Y 0.05fF
C4 w_n6_n6# Y 0.15fF
C5 gnd a_7_n61# 0.45fF
C6 B Y 0.24fF
C7 w_n6_n6# A 0.06fF
C8 B a_7_n61# 0.05fF
C9 vdd Y 1.60fF
C10 w_n6_n6# B 0.06fF

.tran 1n 20n 

.measure tran t_in WHEN v(B)=0.5*SUPPLY CROSS=3
.measure tran t_out WHEN v(Y)=0.5*SUPPLY CROSS=1
.measure tran t_delay PARAM='t_out-t_in'

.control
    set hcopypscolor = 1
    set color0=beige
    set color1=black
    set color2=blue
    set color3=darkgreen
    set color4=darkred
    set color5=darkviolet
    set color6=darkorange

    run
    plot v(A)+4 v(B)+2 v(Y)
.endc