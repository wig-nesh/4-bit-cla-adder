* SPICE3 file created from nor_cmos.ext - technology: scmos

.option scale=0.09u

M1000 a_7_0# A vdd w_n6_n6# pfet w=100 l=2
+  ad=1000 pd=420 as=500 ps=210
M1001 Y B a_7_0# w_n6_n6# pfet w=100 l=2
+  ad=500 pd=210 as=0 ps=0
M1002 Y A gnd Gnd nfet w=20 l=2
+  ad=200 pd=100 as=200 ps=100
M1003 Y B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 A Y 0.05fF
C1 a_7_0# Y 1.03fF
C2 a_7_0# B 0.02fF
C3 a_7_0# vdd 1.03fF
C4 Y gnd 0.71fF
C5 Y w_n6_n6# 0.12fF
C6 B w_n6_n6# 0.06fF
C7 A gnd 0.05fF
C8 A w_n6_n6# 0.06fF
C9 w_n6_n6# vdd 0.12fF
C10 Y B 0.24fF
C11 a_7_0# w_n6_n6# 0.22fF
C12 gnd Gnd 0.15fF
C13 Y Gnd 0.15fF
C14 a_7_0# Gnd 0.00fF
C15 vdd Gnd 0.01fF
C16 B Gnd 0.17fF
C17 A Gnd 0.17fF
C18 w_n6_n6# Gnd 4.50fF
