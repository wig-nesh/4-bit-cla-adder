.include ../../../../tech_files/TSMC_180nm.txt

.param SUPPLY=1.8
.global gnd vdd


VDD vdd gnd SUPPLY
vinA A gnd PULSE(0 SUPPLY 10ns 1ps 1ps 10ns 20ns)

.option scale=0.09u

M1000 OUT IN vdd w_0_0# CMOSP w=50 l=2
+  ad=250 pd=110 as=250 ps=110
M1001 OUT IN gnd Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=100 ps=50
C1 OUT w_0_0# 0.07fF
C2 vdd IN 0.02fF
C3 gnd OUT 0.24fF
C4 OUT IN 0.05fF
C5 IN w_0_0# 0.06fF
C6 vdd OUT 0.55fF
C7 vdd w_0_0# 0.10fF
C8 gnd Gnd 0.12fF
C9 OUT Gnd 0.07fF
C10 vdd Gnd 0.07fF
C11 IN Gnd 0.13fF
C12 w_0_0# Gnd 1.49fF

.tran 1n 20n 

.measure tran t_in WHEN v(A)=0.5*SUPPLY CROSS=1
.measure tran t_out WHEN v(Y)=0.5*SUPPLY CROSS=1
.measure tran t_delay PARAM='t_out-t_in'

.control
    set hcopypscolor = 1
    set color0=beige
    set color1=black
    set color2=blue
    set color3=darkgreen
    set color4=darkred
    set color5=darkviolet
    set color6=darkorange

    run
    plot v(A)+2 v(Y)
.endc