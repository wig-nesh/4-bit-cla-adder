* SPICE3 file created from nand_5_cmos.ext - technology: scmos

.option scale=0.09u

M1000 a_39_n62# C a_23_n62# Gnd nfet w=20 l=2
+  ad=200 pd=100 as=200 ps=100
M1001 a_7_0# A vdd w_n6_n6# pfet w=50 l=2
+  ad=1000 pd=440 as=1250 ps=550
M1002 a_7_0# C vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_7_0# B vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_55_n62# D a_39_n62# Gnd nfet w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1005 Y E a_55_n62# Gnd nfet w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1006 Y E vdd w_n6_n6# pfet w=50 l=2
+  ad=250 pd=110 as=0 ps=0
M1007 a_7_n62# A gnd Gnd nfet w=20 l=2
+  ad=200 pd=100 as=100 ps=50
M1008 a_7_0# D vdd w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_23_n62# B a_7_n62# Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 C B 0.49fF
C1 D A 0.08fF
C2 w_n6_n6# Y 0.07fF
C3 A B 0.27fF
C4 D w_n6_n6# 0.06fF
C5 w_n6_n6# B 0.06fF
C6 Y a_55_n62# 0.21fF
C7 a_23_n62# a_39_n62# 0.21fF
C8 Y E 0.05fF
C9 a_7_0# vdd 4.35fF
C10 C a_7_0# 0.08fF
C11 gnd Y 0.03fF
C12 D E 0.93fF
C13 a_7_0# A 0.05fF
C14 E B 0.08fF
C15 vdd A 0.02fF
C16 a_39_n62# a_55_n62# 0.21fF
C17 C A 0.08fF
C18 a_39_n62# E 0.16fF
C19 w_n6_n6# a_7_0# 0.29fF
C20 w_n6_n6# vdd 0.45fF
C21 a_39_n62# gnd 0.07fF
C22 a_23_n62# a_7_n62# 0.21fF
C23 C w_n6_n6# 0.06fF
C24 w_n6_n6# A 0.06fF
C25 a_7_0# E 0.05fF
C26 C E 0.08fF
C27 a_7_n62# E 0.16fF
C28 E A 0.08fF
C29 D B 0.08fF
C30 gnd a_7_n62# 0.27fF
C31 a_23_n62# E 0.16fF
C32 w_n6_n6# E 0.06fF
C33 a_23_n62# gnd 0.07fF
C34 a_7_0# Y 0.05fF
C35 Y vdd 0.55fF
C36 E a_55_n62# 0.16fF
C37 D a_7_0# 0.08fF
C38 gnd a_55_n62# 0.07fF
C39 a_7_0# B 0.26fF
C40 C D 0.71fF
C41 gnd E 0.05fF
