.include ../../../../tech_files/TSMC_180nm.txt

.param SUPPLY=1.8
.global gnd vdd

VDD vdd gnd SUPPLY
vinA A gnd PULSE(0 SUPPLY  10ns 1ps 1ps  10ns 20ns)
vinB B gnd PULSE(0 SUPPLY   5ns 1ps 1ps   5ns 10ns)
vinC C gnd PULSE(0 SUPPLY 2.5ns 1ps 1ps 2.5ns  5ns)

.option scale=0.09u

M1000 Y A vdd w_n6_n6# CMOSP w=50 l=2
+  ad=750 pd=330 as=750 ps=330
M1001 Y C vdd w_n6_n6# CMOSP w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 Y B vdd w_n6_n6# CMOSP w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_7_n48# A gnd Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=100 ps=50
M1004 a_23_n48# B a_7_n48# Gnd CMOSN w=20 l=2
+  ad=200 pd=100 as=0 ps=0
M1005 Y C a_23_n48# Gnd CMOSN w=20 l=2
+  ad=100 pd=50 as=0 ps=0
C0 A B 0.27fF
C1 Y vdd 2.72fF
C2 C B 0.49fF
C3 w_n6_n6# B 0.06fF
C4 gnd Y 0.03fF
C5 a_23_n48# Y 0.21fF
C6 a_7_n48# gnd 0.27fF
C7 a_23_n48# gnd 0.07fF
C8 vdd A 0.02fF
C9 a_23_n48# a_7_n48# 0.21fF
C10 w_n6_n6# vdd 0.27fF
C11 Y A 0.05fF
C12 Y C 0.13fF
C13 w_n6_n6# Y 0.22fF
C14 gnd C 0.05fF
C15 a_7_n48# C 0.16fF
C16 a_23_n48# C 0.16fF
C17 Y B 0.26fF
C18 A C 0.08fF
C19 w_n6_n6# A 0.06fF
C20 w_n6_n6# C 0.06fF

.tran 1n 20n 

.control
    set hcopypscolor = 1
    set color0=beige
    set color1=black
    set color2=blue
    set color3=darkgreen
    set color4=darkred
    set color5=darkviolet
    set color6=darkorange

    run
    plot v(A)+4 v(B)+2 v(C) v(Y)-2
.endc