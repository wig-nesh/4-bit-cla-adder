magic
tech scmos
timestamp 1731226851
<< nwell >>
rect 0 0 24 62
<< ntransistor >>
rect 11 -28 13 -8
<< ptransistor >>
rect 11 6 13 56
<< ndiffusion >>
rect 10 -28 11 -8
rect 13 -28 14 -8
<< pdiffusion >>
rect 10 6 11 56
rect 13 6 14 56
<< ndcontact >>
rect 6 -28 10 -8
rect 14 -28 18 -8
<< pdcontact >>
rect 6 6 10 56
rect 14 6 18 56
<< polysilicon >>
rect 11 56 13 59
rect 11 -8 13 6
rect 11 -31 13 -28
<< polycontact >>
rect 7 -5 11 -1
<< metal1 >>
rect 6 56 10 65
rect 3 -5 7 -1
rect 14 -8 18 6
rect 6 -37 10 -28
<< labels >>
rlabel metal1 3 -5 7 -1 1 IN
rlabel metal1 14 -5 18 -1 1 OUT
rlabel metal1 6 61 10 65 5 vdd
rlabel metal1 6 -37 10 -33 1 gnd
<< end >>
