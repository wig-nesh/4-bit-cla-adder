* SPICE3 file created from nor_3_cmos.ext - technology: scmos

.option scale=0.09u

M1000 a_7_0# C vdd w_n6_n6# pfet w=50 l=2
+  ad=500 pd=220 as=250 ps=110
M1001 Y A a_23_0# w_n6_n6# pfet w=50 l=2
+  ad=250 pd=110 as=500 ps=220
M1002 a_23_0# B a_7_0# w_n6_n6# pfet w=50 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 Y C gnd Gnd nfet w=20 l=2
+  ad=300 pd=150 as=300 ps=150
M1004 Y B gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 Y A gnd Gnd nfet w=20 l=2
+  ad=0 pd=0 as=0 ps=0
C0 B C 0.27fF
C1 Y B 0.26fF
C2 B A 0.49fF
C3 w_n6_n6# B 0.06fF
C4 a_7_0# vdd 0.61fF
C5 a_23_0# vdd 0.10fF
C6 a_7_0# a_23_0# 0.52fF
C7 C gnd 0.05fF
C8 Y gnd 1.24fF
C9 Y vdd 0.03fF
C10 A vdd 0.02fF
C11 Y a_23_0# 0.52fF
C12 a_7_0# A 0.05fF
C13 a_23_0# A 0.05fF
C14 w_n6_n6# vdd 0.16fF
C15 a_7_0# w_n6_n6# 0.12fF
C16 a_23_0# w_n6_n6# 0.12fF
C17 Y C 0.05fF
C18 C A 0.08fF
C19 w_n6_n6# C 0.06fF
C20 Y A 0.13fF
C21 Y w_n6_n6# 0.07fF
C22 w_n6_n6# A 0.06fF
C23 gnd Gnd 0.32fF
C24 Y Gnd 0.28fF
C25 a_23_0# Gnd 0.00fF
C26 a_7_0# Gnd 0.00fF
C27 vdd Gnd 0.12fF
C28 A Gnd 0.32fF
C29 B Gnd 0.28fF
C30 C Gnd 0.23fF
C31 w_n6_n6# Gnd 3.55fF
