magic
tech scmos
timestamp 1731241506
<< nwell >>
rect -6 -6 82 256
<< ntransistor >>
rect 5 -41 7 -21
rect 21 -41 23 -21
rect 37 -41 39 -21
rect 53 -41 55 -21
rect 69 -41 71 -21
<< ptransistor >>
rect 5 0 7 250
rect 21 0 23 250
rect 37 0 39 250
rect 53 0 55 250
rect 69 0 71 250
<< ndiffusion >>
rect 4 -41 5 -21
rect 7 -41 8 -21
rect 20 -41 21 -21
rect 23 -41 24 -21
rect 36 -41 37 -21
rect 39 -41 40 -21
rect 52 -41 53 -21
rect 55 -41 56 -21
rect 68 -41 69 -21
rect 71 -41 72 -21
<< pdiffusion >>
rect 4 0 5 250
rect 7 0 8 250
rect 20 0 21 250
rect 23 0 24 250
rect 36 0 37 250
rect 39 0 40 250
rect 52 0 53 250
rect 55 0 56 250
rect 68 0 69 250
rect 71 0 72 250
<< ndcontact >>
rect 0 -41 4 -21
rect 8 -41 12 -21
rect 16 -41 20 -21
rect 24 -41 28 -21
rect 32 -41 36 -21
rect 40 -41 44 -21
rect 48 -41 52 -21
rect 56 -41 60 -21
rect 64 -41 68 -21
rect 72 -41 76 -21
<< pdcontact >>
rect 0 0 4 250
rect 8 0 12 250
rect 16 0 20 250
rect 24 0 28 250
rect 32 0 36 250
rect 40 0 44 250
rect 48 0 52 250
rect 56 0 60 250
rect 64 0 68 250
rect 72 0 76 250
<< polysilicon >>
rect 5 250 7 253
rect 21 250 23 253
rect 37 250 39 253
rect 53 250 55 253
rect 69 250 71 253
rect 5 -21 7 0
rect 21 -21 23 0
rect 37 -21 39 0
rect 53 -21 55 0
rect 69 -21 71 0
rect 5 -44 7 -41
rect 21 -44 23 -41
rect 37 -44 39 -41
rect 53 -44 55 -41
rect 69 -44 71 -41
<< polycontact >>
rect 1 -18 5 -14
rect 17 -11 21 -7
rect 33 -11 37 -7
rect 49 -11 53 -7
rect 65 -11 69 -7
<< metal1 >>
rect 0 250 4 259
rect 12 246 16 250
rect 28 246 32 250
rect 44 246 48 250
rect 60 246 64 250
rect 13 -11 17 -7
rect 29 -11 33 -7
rect 45 -11 49 -7
rect 61 -11 65 -7
rect 72 -14 76 0
rect -3 -18 1 -14
rect 8 -18 76 -14
rect 8 -21 12 -18
rect 24 -21 28 -18
rect 40 -21 44 -18
rect 56 -21 60 -18
rect 72 -21 76 -18
rect 0 -46 4 -41
rect 16 -46 20 -41
rect 32 -46 36 -41
rect 48 -46 52 -41
rect 64 -46 68 -41
rect 0 -50 68 -46
<< labels >>
rlabel metal1 61 -11 65 -7 1 E
rlabel metal1 45 -11 49 -7 1 D
rlabel metal1 29 -11 33 -7 1 C
rlabel metal1 13 -11 17 -7 1 B
rlabel metal1 10 -50 14 -46 1 gnd
rlabel metal1 -3 -18 1 -14 1 A
rlabel metal1 72 -11 76 -7 1 Y
rlabel metal1 0 255 4 259 5 vdd
<< end >>
