.include ../../tech_files/TSMC_180nm.txt
.include ../../ckt_blocks/d_ff/optimized/d_ff_optimized.cir
.include ../../ckt_blocks/pg_gen/optimized/pg_gen_optimized.cir
.include ../../ckt_blocks/cla_gen/cmos/cla_gen_cmos.cir
.include ../../ckt_blocks/sum_gen/optimized/sum_gen_optimized.cir

.param SUPPLY=1.8
.param LAMBDA=0.09u
.param width_N={20*LAMBDA}
.param width_P={2.5*width_N}
.param length={2*LAMBDA}
.global gnd vdd

VDD vdd gnd SUPPLY
vinClk clk gnd PULSE(0 SUPPLY 2ns 1ps 1ps 2ns 4ns)
vinA3 A3 gnd PWL(1.99ns 0V 2ns SUPPLY 10.99ns SUPPLY 11ns 0)
vinA2 A2 gnd PWL(1.99ns 0V 2ns SUPPLY 10.99ns SUPPLY 11ns 0)
vinA1 A1 gnd PWL(1.99ns 0V 2ns SUPPLY 10.99ns SUPPLY 11ns 0)
vinA0 A0 gnd PWL(1.99ns 0V 2ns SUPPLY 10.99ns SUPPLY 11ns 0)
vinB3 B3 gnd PWL(1.99ns 0V 2ns SUPPLY 10.99ns SUPPLY 11ns 0)
vinB2 B2 gnd PWL(1.99ns 0V 2ns SUPPLY 10.99ns SUPPLY 11ns 0)
vinB1 B1 gnd PWL(1.99ns 0V 2ns SUPPLY 10.99ns SUPPLY 11ns 0)
vinB0 B0 gnd PWL(1.99ns 0V 2ns SUPPLY 10.99ns SUPPLY 11ns 0)
vinC0 C0 gnd PWL(1.99ns 0V 2ns SUPPLY 10.99ns SUPPLY 11ns 0)

Xdffa3 A3 clk Q3a d_ff_optimized
Xdffa2 A2 clk Q2a d_ff_optimized
Xdffa1 A1 clk Q1a d_ff_optimized
Xdffa0 A0 clk Q0a d_ff_optimized
Xdffb3 B3 clk Q3b d_ff_optimized
Xdffb2 B2 clk Q2b d_ff_optimized
Xdffb1 B1 clk Q1b d_ff_optimized
Xdffb0 B0 clk Q0b d_ff_optimized
Xdffc0 C0 clk Qc0 d_ff_optimized

Xpg  Q3a Q2a Q1a Q0a Q3b Q2b Q1b Q0b P3 P2 P1 P0 G3 G2 G1 G0 pg_gen_optimized
Xcla Qc0  G0  P0  P1  G1  P2  G2  P3 G3 C1 C2 C3 C4 cla_gen_cmos
Xsum  P3  P2  P1  P0  C3  C2  C1  C0 S3 S2 S1 S0 sum_gen_optimized

Xdffs3 S3 clk Q3s d_ff_optimized
Xdffs2 S2 clk Q2s d_ff_optimized
Xdffs1 S1 clk Q1s d_ff_optimized
Xdffs0 S0 clk Q0s d_ff_optimized
Xdffco C4 clk Qco d_ff_optimized

.tran 1n 20n 

.measure tran delay_S3_r TRIG V(A3) VAL=0.5*SUPPLY RISE=1 TARG V(S3) VAL=0.5*SUPPLY RISE=1
.measure tran delay_S2_r TRIG V(A2) VAL=0.5*SUPPLY RISE=1 TARG V(S2) VAL=0.5*SUPPLY RISE=1
.measure tran delay_S1_r TRIG V(A1) VAL=0.5*SUPPLY RISE=1 TARG V(S1) VAL=0.5*SUPPLY RISE=1
.measure tran delay_S0_r TRIG V(A0) VAL=0.5*SUPPLY RISE=1 TARG V(S0) VAL=0.5*SUPPLY RISE=1
.measure tran delay_C4_r TRIG V(C0) VAL=0.5*SUPPLY RISE=1 TARG V(C4) VAL=0.5*SUPPLY RISE=1
.measure tran delay_S3_f TRIG V(A3) VAL=0.5*SUPPLY FALL=1 TARG V(S3) VAL=0.5*SUPPLY FALL=1
.measure tran delay_S2_f TRIG V(A2) VAL=0.5*SUPPLY FALL=1 TARG V(S2) VAL=0.5*SUPPLY FALL=1
.measure tran delay_S1_f TRIG V(A1) VAL=0.5*SUPPLY FALL=1 TARG V(S1) VAL=0.5*SUPPLY FALL=1
.measure tran delay_S0_f TRIG V(A0) VAL=0.5*SUPPLY FALL=1 TARG V(S0) VAL=0.5*SUPPLY FALL=1
.measure tran delay_C4_f TRIG V(C0) VAL=0.5*SUPPLY FALL=1 TARG V(C4) VAL=0.5*SUPPLY FALL=1


.control
    set hcopypscolor = 1
    set color0=beige
    set color1=black
    set color2=blue
    set color3=darkgreen
    set color4=darkgreen
    set color5=darkgreen
    set color6=darkgreen
    set color7=darkred
    set color8=darkred
    set color9=darkred
    set color10=darkred
    set color11=darkviolet
    set color12=darkorange
    set color13=yellow
    set color14=darkorange
    set color15=yellow
    set color16=darkorange
    set color17=yellow
    set color18=darkorange
    set color19=yellow
    set color20=red
    set color21=red
    * set hcopypscolor = 1
    * set color0=beige
    * set color1=black
    * set color2=blue
    * set color3=darkgreen
    * set color4=darkgreen
    * set color5=darkgreen
    * set color6=darkgreen
    * set color7=darkred
    * set color8=darkred
    * set color9=darkred
    * set color10=darkred
    * set color11=darkviolet
    * set color12=darkorange
    * set color13=darkorange
    * set color14=darkorange
    * set color15=darkorange
    * set color16=red
    
    run
    * plot v(clk)+28 v(A3)+26 v(A2)+24 v(A1)+22 v(A0)+20 v(B3)+18 v(B2)+16 v(B1)+14 v(B0)+12 v(C0)+10 v(Q3s)+8 v(S3)+8 v(Q2s)+6 v(S2)+6 v(Q1s)+4 v(S1)+4 v(Q0s)+2 v(S0)+2 v(Qco) v(C4)
    plot v(clk)+28 v(A3)+26 v(A2)+24 v(A1)+22 v(A0)+20 v(B3)+18 v(B2)+16 v(B1)+14 v(B0)+12 v(C0)+10 v(Q3s)+8 v(Q2s)+6 v(Q1s)+4 v(Q0s)+2 v(Qco)
    * plot v(clk)+28 v(A3)+26 v(A2)+24 v(A1)+22 v(A0)+20 v(B3)+18 v(B2)+16 v(B1)+14 v(B0)+12 v(C0)+10 v(Q3s)+8 v(Q2s)+6 v(Q1s)+4 v(Q0s)+2 v(Qco)
    set curplottitle="2023102019"
    hardcopy full_optimized_tran.eps v(clk)+28 v(A3)+26 v(A2)+24 v(A1)+22 v(A0)+20 v(B3)+18 v(B2)+16 v(B1)+14 v(B0)+12 v(C0)+10 v(Q3s)+8 v(Q2s)+6 v(Q1s)+4 v(Q0s)+2 v(Qco)
.endc   